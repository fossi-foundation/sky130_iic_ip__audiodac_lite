magic
tech sky130A
magscale 1 2
timestamp 1645182741
<< nwell >>
rect 222554 108114 222874 108366
rect 222542 108094 222874 108114
rect 222542 107358 222832 108094
rect 222562 106124 222830 107358
rect 222562 104140 222828 106124
rect 222548 103558 222870 104140
rect 222548 103536 223082 103558
rect 222572 103530 223082 103536
rect 222550 84836 222642 84838
rect 222550 84818 223068 84836
rect 222550 84808 222854 84818
rect 222516 81242 222854 84808
rect 222522 80218 222854 81242
rect 222522 80046 222918 80218
rect 222456 80000 222990 80046
<< locali >>
rect 220138 90632 220278 91300
rect 222318 91280 222466 91302
rect 220142 80304 220276 90632
rect 222318 80342 222470 91280
rect 220142 80298 220294 80304
rect 220144 80292 220294 80298
rect 222318 80292 222472 80342
<< metal1 >>
rect 220278 103206 220288 105232
rect 222362 103206 222372 105232
rect 223364 101278 223370 101386
rect 223478 101278 223484 101386
rect 222719 98784 222986 98974
rect 220314 96928 220324 97048
rect 222322 96928 222332 97048
rect 222719 95727 222909 98784
rect 222719 95537 223407 95727
rect 220022 92929 220124 95196
rect 223217 93773 223407 95537
rect 223217 93583 223681 93773
rect 224370 93604 224808 93764
rect 224648 92132 224808 93604
rect 223950 91972 224808 92132
rect 223950 91956 224110 91972
rect 222796 91796 224110 91956
rect 220296 91346 220306 91440
rect 222306 91346 222316 91440
rect 222796 89236 222956 91796
rect 223364 86934 223370 87042
rect 223478 86934 223484 87042
rect 220250 83680 220260 85652
rect 222356 83680 222366 85652
<< via1 >>
rect 220288 103206 222362 105232
rect 223370 101278 223478 101386
rect 220324 96928 222322 97048
rect 220306 91346 222306 91440
rect 223370 86934 223478 87042
rect 220260 83680 222356 85652
<< metal2 >>
rect 220288 105232 222362 105242
rect 220288 103196 222362 103206
rect 223370 101386 223478 101392
rect 223361 101278 223370 101386
rect 223478 101278 223487 101386
rect 223370 101272 223478 101278
rect 225000 99890 225100 99899
rect 225000 99721 225100 99730
rect 220320 97048 225042 97468
rect 220320 96928 220324 97048
rect 222322 96928 225042 97048
rect 220320 96852 225042 96928
rect 222567 96057 222631 96091
rect 222567 96056 222742 96057
rect 222567 95975 222852 96056
rect 222567 95971 222631 95975
rect 222742 95917 222852 95975
rect 224595 95960 224765 95969
rect 223907 95917 223989 95960
rect 222742 95836 223989 95917
rect 222852 95835 223989 95836
rect 220994 95701 221003 95799
rect 221101 95701 221110 95799
rect 222145 95789 222243 95798
rect 223907 95790 223989 95835
rect 224221 95790 224595 95960
rect 224595 95781 224765 95790
rect 222145 95682 222243 95691
rect 223591 92536 223855 92576
rect 223116 92412 225008 92536
rect 223116 92286 223240 92412
rect 223591 92406 223855 92412
rect 220565 92161 220705 92285
rect 222686 92162 223240 92286
rect 224884 91540 225008 92412
rect 220298 91440 225066 91540
rect 220298 91346 220306 91440
rect 222306 91346 225066 91440
rect 220298 91152 225066 91346
rect 223370 87042 223478 87048
rect 223361 86934 223370 87042
rect 223478 86934 223487 87042
rect 223370 86928 223478 86934
rect 220260 85652 222356 85662
rect 220260 83670 222356 83680
<< via2 >>
rect 220288 103206 222362 105232
rect 223370 101278 223478 101386
rect 221003 95701 221101 95799
rect 224595 95790 224765 95960
rect 222145 95691 222243 95789
rect 223370 86934 223478 87042
rect 220260 83680 222356 85652
<< metal3 >>
rect 220288 105237 228486 105260
rect 220278 105232 228486 105237
rect 220278 103206 220288 105232
rect 222362 103206 228486 105232
rect 220278 103201 222372 103206
rect 228720 101846 232044 106696
rect 223365 101386 223483 101391
rect 222830 101278 223370 101386
rect 223478 101278 223483 101386
rect 222830 96150 222938 101278
rect 223365 101273 223483 101278
rect 228720 101046 232052 101846
rect 232502 101092 234338 102848
rect 220998 96042 222938 96150
rect 225454 99650 228538 99712
rect 220998 95799 221106 96042
rect 225454 95966 225498 99650
rect 220998 95701 221003 95799
rect 221101 95701 221106 95799
rect 224584 95960 225498 95966
rect 220998 95688 221106 95701
rect 222140 95789 223186 95794
rect 222140 95691 222145 95789
rect 222243 95691 223186 95789
rect 224584 95790 224595 95960
rect 224765 95790 225498 95960
rect 224584 95780 225498 95790
rect 222140 95686 223186 95691
rect 220091 92509 222771 92589
rect 220091 92329 220381 92409
rect 223078 92006 223186 95686
rect 222832 91898 223186 92006
rect 225454 95100 225498 95780
rect 228460 95100 228538 99650
rect 228728 96610 232052 101046
rect 222832 87042 222940 91898
rect 223365 87042 223483 87047
rect 222832 86934 223370 87042
rect 223478 86934 223483 87042
rect 223365 86929 223483 86934
rect 225454 86526 228538 95100
rect 228724 96196 232052 96610
rect 228724 93336 232048 96196
rect 228724 91358 228854 93336
rect 220250 85652 228470 85662
rect 220250 83680 220260 85652
rect 222356 83680 228470 85652
rect 220250 83676 228470 83680
rect 220250 83675 222366 83676
rect 228738 81868 228854 91358
rect 231886 92020 232048 93336
rect 231886 81868 232062 92020
rect 232502 85518 234338 87274
rect 228738 81720 232062 81868
<< via3 >>
rect 225498 95100 228460 99650
rect 228854 81868 231886 93336
<< metal4 >>
rect 220092 106932 234472 108248
rect 220092 99650 234472 105846
rect 220092 95100 225498 99650
rect 228460 95100 234472 99650
rect 220092 95044 234472 95100
rect 220092 93336 234472 93464
rect 220092 89374 228854 93336
rect 231886 89374 234472 93336
rect 234448 88214 234472 89374
rect 220092 81868 228854 88214
rect 231886 81868 234472 88214
rect 220092 80260 234472 81868
<< via4 >>
rect 220070 105846 234740 106932
rect 220054 88214 228854 89374
rect 228854 88214 231886 89374
rect 231886 88214 234448 89374
<< metal5 >>
rect 220046 106932 234764 106956
rect 220046 105846 220070 106932
rect 234740 105846 234764 106932
rect 220046 105822 234764 105846
rect 220030 89374 234472 89398
rect 220030 88214 220054 89374
rect 234448 88214 234472 89374
rect 220030 88190 234472 88214
use audiodac_drv_half  audiodac_drv_half_0
timestamp 1644660203
transform 1 0 228698 0 1 115642
box -5906 -21361 6044 -7276
use audiodac_drv_half  audiodac_drv_half_1
timestamp 1644660203
transform 1 0 228698 0 -1 72724
box -5906 -21361 6044 -7276
use audiodac_drv_latch  audiodac_drv_latch_0
timestamp 1644659262
transform 1 0 221501 0 1 119112
box 1834 -27002 3224 -22840
use audiodac_drv_ls  audiodac_drv_ls_0
timestamp 1644660372
transform 1 0 223749 0 1 111945
box -3728 -20005 -570 -15559
use jku_logo  jku_logo_0
timestamp 1645179649
transform 1 0 -46 0 1 1960
box 338 0 234514 75214
use sky130_fd_pr__pfet_g5v0d10v5_VDASXE  sky130_fd_pr__pfet_g5v0d10v5_VDASXE_0  paramcells
timestamp 1644523392
transform 1 0 221326 0 1 102589
box -1258 -5797 1258 5797
use sky130_fd_pr__pfet_g5v0d10v5_VDASXE  sky130_fd_pr__pfet_g5v0d10v5_VDASXE_1
timestamp 1644523392
transform 1 0 221306 0 1 85797
box -1258 -5797 1258 5797
<< labels >>
rlabel metal3 220091 92509 222771 92589 1 in_n
port 2 n signal input
rlabel metal3 220091 92329 220381 92409 1 in_p
port 1 n signal input
rlabel metal3 232502 85518 234338 87274 1 out_p
port 3 n signal output
rlabel metal3 232502 101092 234338 102848 1 out_n
port 4 n signal output
rlabel metal3 228738 81720 232062 92020 1 vss
port 7 n ground input
rlabel metal3 225454 86526 228538 99712 1 vdd
port 5 n power input
rlabel metal1 220022 92929 220124 95196 1 in_hi
port 6 n signal input
<< end >>
