magic
tech sky130A
timestamp 1644523392
<< pwell >>
rect -257 -379 257 379
<< mvnmos >>
rect -143 -250 -93 250
rect -64 -250 -14 250
rect 15 -250 65 250
rect 94 -250 144 250
<< mvndiff >>
rect -172 244 -143 250
rect -172 -244 -166 244
rect -149 -244 -143 244
rect -172 -250 -143 -244
rect -93 244 -64 250
rect -93 -244 -87 244
rect -70 -244 -64 244
rect -93 -250 -64 -244
rect -14 244 15 250
rect -14 -244 -8 244
rect 9 -244 15 244
rect -14 -250 15 -244
rect 65 244 94 250
rect 65 -244 71 244
rect 88 -244 94 244
rect 65 -250 94 -244
rect 144 244 173 250
rect 144 -244 150 244
rect 167 -244 173 244
rect 144 -250 173 -244
<< mvndiffc >>
rect -166 -244 -149 244
rect -87 -244 -70 244
rect -8 -244 9 244
rect 71 -244 88 244
rect 150 -244 167 244
<< mvpsubdiff >>
rect -239 355 239 361
rect -239 338 -185 355
rect 185 338 239 355
rect -239 332 239 338
rect -239 307 -210 332
rect -239 -307 -233 307
rect -216 -307 -210 307
rect 210 307 239 332
rect -239 -332 -210 -307
rect 210 -307 216 307
rect 233 -307 239 307
rect 210 -332 239 -307
rect -239 -338 239 -332
rect -239 -355 -185 -338
rect 185 -355 239 -338
rect -239 -361 239 -355
<< mvpsubdiffcont >>
rect -185 338 185 355
rect -233 -307 -216 307
rect 216 -307 233 307
rect -185 -355 185 -338
<< poly >>
rect -143 286 -93 294
rect -143 269 -135 286
rect -101 269 -93 286
rect -143 250 -93 269
rect -64 286 -14 294
rect -64 269 -56 286
rect -22 269 -14 286
rect -64 250 -14 269
rect 15 286 65 294
rect 15 269 23 286
rect 57 269 65 286
rect 15 250 65 269
rect 94 286 144 294
rect 94 269 102 286
rect 136 269 144 286
rect 94 250 144 269
rect -143 -269 -93 -250
rect -143 -286 -135 -269
rect -101 -286 -93 -269
rect -143 -294 -93 -286
rect -64 -269 -14 -250
rect -64 -286 -56 -269
rect -22 -286 -14 -269
rect -64 -294 -14 -286
rect 15 -269 65 -250
rect 15 -286 23 -269
rect 57 -286 65 -269
rect 15 -294 65 -286
rect 94 -269 144 -250
rect 94 -286 102 -269
rect 136 -286 144 -269
rect 94 -294 144 -286
<< polycont >>
rect -135 269 -101 286
rect -56 269 -22 286
rect 23 269 57 286
rect 102 269 136 286
rect -135 -286 -101 -269
rect -56 -286 -22 -269
rect 23 -286 57 -269
rect 102 -286 136 -269
<< locali >>
rect -233 338 -185 355
rect 185 338 233 355
rect -233 307 -216 338
rect 216 307 233 338
rect -143 269 -135 286
rect -101 269 -93 286
rect -64 269 -56 286
rect -22 269 -14 286
rect 15 269 23 286
rect 57 269 65 286
rect 94 269 102 286
rect 136 269 144 286
rect -166 244 -149 252
rect -166 -252 -149 -244
rect -87 244 -70 252
rect -87 -252 -70 -244
rect -8 244 9 252
rect -8 -252 9 -244
rect 71 244 88 252
rect 71 -252 88 -244
rect 150 244 167 252
rect 150 -252 167 -244
rect -143 -286 -135 -269
rect -101 -286 -93 -269
rect -64 -286 -56 -269
rect -22 -286 -14 -269
rect 15 -286 23 -269
rect 57 -286 65 -269
rect 94 -286 102 -269
rect 136 -286 144 -269
rect -233 -338 -216 -307
rect 216 -338 233 -307
rect -233 -355 -185 -338
rect 185 -355 233 -338
<< viali >>
rect -135 269 -101 286
rect -56 269 -22 286
rect 23 269 57 286
rect 102 269 136 286
rect -166 -244 -149 244
rect -87 -244 -70 244
rect -8 -244 9 244
rect 71 -244 88 244
rect 150 -244 167 244
rect -135 -286 -101 -269
rect -56 -286 -22 -269
rect 23 -286 57 -269
rect 102 -286 136 -269
<< metal1 >>
rect -141 286 -95 289
rect -141 269 -135 286
rect -101 269 -95 286
rect -141 266 -95 269
rect -62 286 -16 289
rect -62 269 -56 286
rect -22 269 -16 286
rect -62 266 -16 269
rect 17 286 63 289
rect 17 269 23 286
rect 57 269 63 286
rect 17 266 63 269
rect 96 286 142 289
rect 96 269 102 286
rect 136 269 142 286
rect 96 266 142 269
rect -169 244 -146 250
rect -169 -244 -166 244
rect -149 -244 -146 244
rect -169 -250 -146 -244
rect -90 244 -67 250
rect -90 -244 -87 244
rect -70 -244 -67 244
rect -90 -250 -67 -244
rect -11 244 12 250
rect -11 -244 -8 244
rect 9 -244 12 244
rect -11 -250 12 -244
rect 68 244 91 250
rect 68 -244 71 244
rect 88 -244 91 244
rect 68 -250 91 -244
rect 147 244 170 250
rect 147 -244 150 244
rect 167 -244 170 244
rect 147 -250 170 -244
rect -141 -269 -95 -266
rect -141 -286 -135 -269
rect -101 -286 -95 -269
rect -141 -289 -95 -286
rect -62 -269 -16 -266
rect -62 -286 -56 -269
rect -22 -286 -16 -269
rect -62 -289 -16 -286
rect 17 -269 63 -266
rect 17 -286 23 -269
rect 57 -286 63 -269
rect 17 -289 63 -286
rect 96 -269 142 -266
rect 96 -286 102 -269
rect 136 -286 142 -269
rect 96 -289 142 -286
<< properties >>
string FIXED_BBOX -225 -346 225 346
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 5 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
