magic
tech sky130A
timestamp 1644523392
<< pwell >>
rect -494 -629 494 629
<< mvnmos >>
rect -380 -500 -330 500
rect -301 -500 -251 500
rect -222 -500 -172 500
rect -143 -500 -93 500
rect -64 -500 -14 500
rect 15 -500 65 500
rect 94 -500 144 500
rect 173 -500 223 500
rect 252 -500 302 500
rect 331 -500 381 500
<< mvndiff >>
rect -409 494 -380 500
rect -409 -494 -403 494
rect -386 -494 -380 494
rect -409 -500 -380 -494
rect -330 494 -301 500
rect -330 -494 -324 494
rect -307 -494 -301 494
rect -330 -500 -301 -494
rect -251 494 -222 500
rect -251 -494 -245 494
rect -228 -494 -222 494
rect -251 -500 -222 -494
rect -172 494 -143 500
rect -172 -494 -166 494
rect -149 -494 -143 494
rect -172 -500 -143 -494
rect -93 494 -64 500
rect -93 -494 -87 494
rect -70 -494 -64 494
rect -93 -500 -64 -494
rect -14 494 15 500
rect -14 -494 -8 494
rect 9 -494 15 494
rect -14 -500 15 -494
rect 65 494 94 500
rect 65 -494 71 494
rect 88 -494 94 494
rect 65 -500 94 -494
rect 144 494 173 500
rect 144 -494 150 494
rect 167 -494 173 494
rect 144 -500 173 -494
rect 223 494 252 500
rect 223 -494 229 494
rect 246 -494 252 494
rect 223 -500 252 -494
rect 302 494 331 500
rect 302 -494 308 494
rect 325 -494 331 494
rect 302 -500 331 -494
rect 381 494 410 500
rect 381 -494 387 494
rect 404 -494 410 494
rect 381 -500 410 -494
<< mvndiffc >>
rect -403 -494 -386 494
rect -324 -494 -307 494
rect -245 -494 -228 494
rect -166 -494 -149 494
rect -87 -494 -70 494
rect -8 -494 9 494
rect 71 -494 88 494
rect 150 -494 167 494
rect 229 -494 246 494
rect 308 -494 325 494
rect 387 -494 404 494
<< mvpsubdiff >>
rect -476 605 476 611
rect -476 588 -422 605
rect 422 588 476 605
rect -476 582 476 588
rect -476 557 -447 582
rect -476 -557 -470 557
rect -453 -557 -447 557
rect 447 557 476 582
rect -476 -582 -447 -557
rect 447 -557 453 557
rect 470 -557 476 557
rect 447 -582 476 -557
rect -476 -588 476 -582
rect -476 -605 -422 -588
rect 422 -605 476 -588
rect -476 -611 476 -605
<< mvpsubdiffcont >>
rect -422 588 422 605
rect -470 -557 -453 557
rect 453 -557 470 557
rect -422 -605 422 -588
<< poly >>
rect -380 536 -330 544
rect -380 519 -372 536
rect -338 519 -330 536
rect -380 500 -330 519
rect -301 536 -251 544
rect -301 519 -293 536
rect -259 519 -251 536
rect -301 500 -251 519
rect -222 536 -172 544
rect -222 519 -214 536
rect -180 519 -172 536
rect -222 500 -172 519
rect -143 536 -93 544
rect -143 519 -135 536
rect -101 519 -93 536
rect -143 500 -93 519
rect -64 536 -14 544
rect -64 519 -56 536
rect -22 519 -14 536
rect -64 500 -14 519
rect 15 536 65 544
rect 15 519 23 536
rect 57 519 65 536
rect 15 500 65 519
rect 94 536 144 544
rect 94 519 102 536
rect 136 519 144 536
rect 94 500 144 519
rect 173 536 223 544
rect 173 519 181 536
rect 215 519 223 536
rect 173 500 223 519
rect 252 536 302 544
rect 252 519 260 536
rect 294 519 302 536
rect 252 500 302 519
rect 331 536 381 544
rect 331 519 339 536
rect 373 519 381 536
rect 331 500 381 519
rect -380 -519 -330 -500
rect -380 -536 -372 -519
rect -338 -536 -330 -519
rect -380 -544 -330 -536
rect -301 -519 -251 -500
rect -301 -536 -293 -519
rect -259 -536 -251 -519
rect -301 -544 -251 -536
rect -222 -519 -172 -500
rect -222 -536 -214 -519
rect -180 -536 -172 -519
rect -222 -544 -172 -536
rect -143 -519 -93 -500
rect -143 -536 -135 -519
rect -101 -536 -93 -519
rect -143 -544 -93 -536
rect -64 -519 -14 -500
rect -64 -536 -56 -519
rect -22 -536 -14 -519
rect -64 -544 -14 -536
rect 15 -519 65 -500
rect 15 -536 23 -519
rect 57 -536 65 -519
rect 15 -544 65 -536
rect 94 -519 144 -500
rect 94 -536 102 -519
rect 136 -536 144 -519
rect 94 -544 144 -536
rect 173 -519 223 -500
rect 173 -536 181 -519
rect 215 -536 223 -519
rect 173 -544 223 -536
rect 252 -519 302 -500
rect 252 -536 260 -519
rect 294 -536 302 -519
rect 252 -544 302 -536
rect 331 -519 381 -500
rect 331 -536 339 -519
rect 373 -536 381 -519
rect 331 -544 381 -536
<< polycont >>
rect -372 519 -338 536
rect -293 519 -259 536
rect -214 519 -180 536
rect -135 519 -101 536
rect -56 519 -22 536
rect 23 519 57 536
rect 102 519 136 536
rect 181 519 215 536
rect 260 519 294 536
rect 339 519 373 536
rect -372 -536 -338 -519
rect -293 -536 -259 -519
rect -214 -536 -180 -519
rect -135 -536 -101 -519
rect -56 -536 -22 -519
rect 23 -536 57 -519
rect 102 -536 136 -519
rect 181 -536 215 -519
rect 260 -536 294 -519
rect 339 -536 373 -519
<< locali >>
rect -470 588 -422 605
rect 422 588 470 605
rect -470 557 -453 588
rect 453 557 470 588
rect -380 519 -372 536
rect -338 519 -330 536
rect -301 519 -293 536
rect -259 519 -251 536
rect -222 519 -214 536
rect -180 519 -172 536
rect -143 519 -135 536
rect -101 519 -93 536
rect -64 519 -56 536
rect -22 519 -14 536
rect 15 519 23 536
rect 57 519 65 536
rect 94 519 102 536
rect 136 519 144 536
rect 173 519 181 536
rect 215 519 223 536
rect 252 519 260 536
rect 294 519 302 536
rect 331 519 339 536
rect 373 519 381 536
rect -403 494 -386 502
rect -403 -502 -386 -494
rect -324 494 -307 502
rect -324 -502 -307 -494
rect -245 494 -228 502
rect -245 -502 -228 -494
rect -166 494 -149 502
rect -166 -502 -149 -494
rect -87 494 -70 502
rect -87 -502 -70 -494
rect -8 494 9 502
rect -8 -502 9 -494
rect 71 494 88 502
rect 71 -502 88 -494
rect 150 494 167 502
rect 150 -502 167 -494
rect 229 494 246 502
rect 229 -502 246 -494
rect 308 494 325 502
rect 308 -502 325 -494
rect 387 494 404 502
rect 387 -502 404 -494
rect -380 -536 -372 -519
rect -338 -536 -330 -519
rect -301 -536 -293 -519
rect -259 -536 -251 -519
rect -222 -536 -214 -519
rect -180 -536 -172 -519
rect -143 -536 -135 -519
rect -101 -536 -93 -519
rect -64 -536 -56 -519
rect -22 -536 -14 -519
rect 15 -536 23 -519
rect 57 -536 65 -519
rect 94 -536 102 -519
rect 136 -536 144 -519
rect 173 -536 181 -519
rect 215 -536 223 -519
rect 252 -536 260 -519
rect 294 -536 302 -519
rect 331 -536 339 -519
rect 373 -536 381 -519
rect -470 -588 -453 -557
rect 453 -588 470 -557
rect -470 -605 -422 -588
rect 422 -605 470 -588
<< viali >>
rect -372 519 -338 536
rect -293 519 -259 536
rect -214 519 -180 536
rect -135 519 -101 536
rect -56 519 -22 536
rect 23 519 57 536
rect 102 519 136 536
rect 181 519 215 536
rect 260 519 294 536
rect 339 519 373 536
rect -403 -494 -386 494
rect -324 -494 -307 494
rect -245 -494 -228 494
rect -166 -494 -149 494
rect -87 -494 -70 494
rect -8 -494 9 494
rect 71 -494 88 494
rect 150 -494 167 494
rect 229 -494 246 494
rect 308 -494 325 494
rect 387 -494 404 494
rect -372 -536 -338 -519
rect -293 -536 -259 -519
rect -214 -536 -180 -519
rect -135 -536 -101 -519
rect -56 -536 -22 -519
rect 23 -536 57 -519
rect 102 -536 136 -519
rect 181 -536 215 -519
rect 260 -536 294 -519
rect 339 -536 373 -519
<< metal1 >>
rect -378 536 -332 539
rect -378 519 -372 536
rect -338 519 -332 536
rect -378 516 -332 519
rect -299 536 -253 539
rect -299 519 -293 536
rect -259 519 -253 536
rect -299 516 -253 519
rect -220 536 -174 539
rect -220 519 -214 536
rect -180 519 -174 536
rect -220 516 -174 519
rect -141 536 -95 539
rect -141 519 -135 536
rect -101 519 -95 536
rect -141 516 -95 519
rect -62 536 -16 539
rect -62 519 -56 536
rect -22 519 -16 536
rect -62 516 -16 519
rect 17 536 63 539
rect 17 519 23 536
rect 57 519 63 536
rect 17 516 63 519
rect 96 536 142 539
rect 96 519 102 536
rect 136 519 142 536
rect 96 516 142 519
rect 175 536 221 539
rect 175 519 181 536
rect 215 519 221 536
rect 175 516 221 519
rect 254 536 300 539
rect 254 519 260 536
rect 294 519 300 536
rect 254 516 300 519
rect 333 536 379 539
rect 333 519 339 536
rect 373 519 379 536
rect 333 516 379 519
rect -406 494 -383 500
rect -406 -494 -403 494
rect -386 -494 -383 494
rect -406 -500 -383 -494
rect -327 494 -304 500
rect -327 -494 -324 494
rect -307 -494 -304 494
rect -327 -500 -304 -494
rect -248 494 -225 500
rect -248 -494 -245 494
rect -228 -494 -225 494
rect -248 -500 -225 -494
rect -169 494 -146 500
rect -169 -494 -166 494
rect -149 -494 -146 494
rect -169 -500 -146 -494
rect -90 494 -67 500
rect -90 -494 -87 494
rect -70 -494 -67 494
rect -90 -500 -67 -494
rect -11 494 12 500
rect -11 -494 -8 494
rect 9 -494 12 494
rect -11 -500 12 -494
rect 68 494 91 500
rect 68 -494 71 494
rect 88 -494 91 494
rect 68 -500 91 -494
rect 147 494 170 500
rect 147 -494 150 494
rect 167 -494 170 494
rect 147 -500 170 -494
rect 226 494 249 500
rect 226 -494 229 494
rect 246 -494 249 494
rect 226 -500 249 -494
rect 305 494 328 500
rect 305 -494 308 494
rect 325 -494 328 494
rect 305 -500 328 -494
rect 384 494 407 500
rect 384 -494 387 494
rect 404 -494 407 494
rect 384 -500 407 -494
rect -378 -519 -332 -516
rect -378 -536 -372 -519
rect -338 -536 -332 -519
rect -378 -539 -332 -536
rect -299 -519 -253 -516
rect -299 -536 -293 -519
rect -259 -536 -253 -519
rect -299 -539 -253 -536
rect -220 -519 -174 -516
rect -220 -536 -214 -519
rect -180 -536 -174 -519
rect -220 -539 -174 -536
rect -141 -519 -95 -516
rect -141 -536 -135 -519
rect -101 -536 -95 -519
rect -141 -539 -95 -536
rect -62 -519 -16 -516
rect -62 -536 -56 -519
rect -22 -536 -16 -519
rect -62 -539 -16 -536
rect 17 -519 63 -516
rect 17 -536 23 -519
rect 57 -536 63 -519
rect 17 -539 63 -536
rect 96 -519 142 -516
rect 96 -536 102 -519
rect 136 -536 142 -519
rect 96 -539 142 -536
rect 175 -519 221 -516
rect 175 -536 181 -519
rect 215 -536 221 -519
rect 175 -539 221 -536
rect 254 -519 300 -516
rect 254 -536 260 -519
rect 294 -536 300 -519
rect 254 -539 300 -536
rect 333 -519 379 -516
rect 333 -536 339 -519
rect 373 -536 379 -519
rect 333 -539 379 -536
<< properties >>
string FIXED_BBOX -462 -596 462 596
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.50 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
