magic
tech sky130A
magscale 1 2
timestamp 1644523201
<< nwell >>
rect -1196 -5719 1196 5719
<< pmos >>
rect -1000 -5500 1000 5500
<< pdiff >>
rect -1058 5488 -1000 5500
rect -1058 -5488 -1046 5488
rect -1012 -5488 -1000 5488
rect -1058 -5500 -1000 -5488
rect 1000 5488 1058 5500
rect 1000 -5488 1012 5488
rect 1046 -5488 1058 5488
rect 1000 -5500 1058 -5488
<< pdiffc >>
rect -1046 -5488 -1012 5488
rect 1012 -5488 1046 5488
<< nsubdiff >>
rect -1160 5649 -1064 5683
rect 1064 5649 1160 5683
rect -1160 5587 -1126 5649
rect 1126 5587 1160 5649
rect -1160 -5649 -1126 -5587
rect 1126 -5649 1160 -5587
rect -1160 -5683 -1064 -5649
rect 1064 -5683 1160 -5649
<< nsubdiffcont >>
rect -1064 5649 1064 5683
rect -1160 -5587 -1126 5587
rect 1126 -5587 1160 5587
rect -1064 -5683 1064 -5649
<< poly >>
rect -1000 5581 1000 5597
rect -1000 5547 -984 5581
rect 984 5547 1000 5581
rect -1000 5500 1000 5547
rect -1000 -5547 1000 -5500
rect -1000 -5581 -984 -5547
rect 984 -5581 1000 -5547
rect -1000 -5597 1000 -5581
<< polycont >>
rect -984 5547 984 5581
rect -984 -5581 984 -5547
<< locali >>
rect -1160 5649 -1064 5683
rect 1064 5649 1160 5683
rect -1160 5587 -1126 5649
rect 1126 5587 1160 5649
rect -1000 5547 -984 5581
rect 984 5547 1000 5581
rect -1046 5488 -1012 5504
rect -1046 -5504 -1012 -5488
rect 1012 5488 1046 5504
rect 1012 -5504 1046 -5488
rect -1000 -5581 -984 -5547
rect 984 -5581 1000 -5547
rect -1160 -5649 -1126 -5587
rect 1126 -5649 1160 -5587
rect -1160 -5683 -1064 -5649
rect 1064 -5683 1160 -5649
<< viali >>
rect -984 5547 984 5581
rect -1046 -5488 -1012 5488
rect 1012 -5488 1046 5488
rect -984 -5581 984 -5547
<< metal1 >>
rect -996 5581 996 5587
rect -996 5547 -984 5581
rect 984 5547 996 5581
rect -996 5541 996 5547
rect -1052 5488 -1006 5500
rect -1052 -5488 -1046 5488
rect -1012 -5488 -1006 5488
rect -1052 -5500 -1006 -5488
rect 1006 5488 1052 5500
rect 1006 -5488 1012 5488
rect 1046 -5488 1052 5488
rect 1006 -5500 1052 -5488
rect -996 -5547 996 -5541
rect -996 -5581 -984 -5547
rect 984 -5581 996 -5547
rect -996 -5587 996 -5581
<< properties >>
string FIXED_BBOX -1143 -5666 1143 5666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 55 l 10 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
