magic
tech sky130A
timestamp 1644523392
<< error_p >>
rect -182 136 -153 139
rect -86 136 -57 139
rect 9 136 38 139
rect 105 136 134 139
rect 201 136 230 139
rect -182 119 -176 136
rect -86 119 -80 136
rect 9 119 15 136
rect 105 119 111 136
rect 201 119 207 136
rect -182 116 -153 119
rect -86 116 -57 119
rect 9 116 38 119
rect 105 116 134 119
rect 201 116 230 119
rect -230 -119 -201 -116
rect -134 -119 -105 -116
rect -38 -119 -9 -116
rect 57 -119 86 -116
rect 153 -119 182 -116
rect -230 -136 -224 -119
rect -134 -136 -128 -119
rect -38 -136 -32 -119
rect 57 -136 63 -119
rect 153 -136 159 -119
rect -230 -139 -201 -136
rect -134 -139 -105 -136
rect -38 -139 -9 -136
rect 57 -139 86 -136
rect 153 -139 182 -136
<< pwell >>
rect -323 -205 323 205
<< nmos >>
rect -223 -100 -208 100
rect -175 -100 -160 100
rect -127 -100 -112 100
rect -79 -100 -64 100
rect -31 -100 -16 100
rect 16 -100 31 100
rect 64 -100 79 100
rect 112 -100 127 100
rect 160 -100 175 100
rect 208 -100 223 100
<< ndiff >>
rect -254 94 -223 100
rect -254 -94 -248 94
rect -231 -94 -223 94
rect -254 -100 -223 -94
rect -208 94 -175 100
rect -208 -94 -200 94
rect -183 -94 -175 94
rect -208 -100 -175 -94
rect -160 94 -127 100
rect -160 -94 -152 94
rect -135 -94 -127 94
rect -160 -100 -127 -94
rect -112 94 -79 100
rect -112 -94 -104 94
rect -87 -94 -79 94
rect -112 -100 -79 -94
rect -64 94 -31 100
rect -64 -94 -56 94
rect -39 -94 -31 94
rect -64 -100 -31 -94
rect -16 94 16 100
rect -16 -94 -8 94
rect 9 -94 16 94
rect -16 -100 16 -94
rect 31 94 64 100
rect 31 -94 39 94
rect 56 -94 64 94
rect 31 -100 64 -94
rect 79 94 112 100
rect 79 -94 87 94
rect 104 -94 112 94
rect 79 -100 112 -94
rect 127 94 160 100
rect 127 -94 135 94
rect 152 -94 160 94
rect 127 -100 160 -94
rect 175 94 208 100
rect 175 -94 183 94
rect 200 -94 208 94
rect 175 -100 208 -94
rect 223 94 254 100
rect 223 -94 231 94
rect 248 -94 254 94
rect 223 -100 254 -94
<< ndiffc >>
rect -248 -94 -231 94
rect -200 -94 -183 94
rect -152 -94 -135 94
rect -104 -94 -87 94
rect -56 -94 -39 94
rect -8 -94 9 94
rect 39 -94 56 94
rect 87 -94 104 94
rect 135 -94 152 94
rect 183 -94 200 94
rect 231 -94 248 94
<< psubdiff >>
rect -305 170 -257 187
rect 257 170 305 187
rect -305 139 -288 170
rect 288 139 305 170
rect -305 -170 -288 -139
rect 288 -170 305 -139
rect -305 -187 -257 -170
rect 257 -187 305 -170
<< psubdiffcont >>
rect -257 170 257 187
rect -305 -139 -288 139
rect 288 -139 305 139
rect -257 -187 257 -170
<< poly >>
rect -184 136 -151 144
rect -184 119 -176 136
rect -159 119 -151 136
rect -223 100 -208 113
rect -184 111 -151 119
rect -88 136 -55 144
rect -88 119 -80 136
rect -63 119 -55 136
rect -175 100 -160 111
rect -127 100 -112 113
rect -88 111 -55 119
rect 7 136 40 144
rect 7 119 15 136
rect 32 119 40 136
rect -79 100 -64 111
rect -31 100 -16 113
rect 7 111 40 119
rect 103 136 136 144
rect 103 119 111 136
rect 128 119 136 136
rect 16 100 31 111
rect 64 100 79 113
rect 103 111 136 119
rect 199 136 232 144
rect 199 119 207 136
rect 224 119 232 136
rect 112 100 127 111
rect 160 100 175 113
rect 199 111 232 119
rect 208 100 223 111
rect -223 -111 -208 -100
rect -232 -119 -199 -111
rect -175 -113 -160 -100
rect -127 -111 -112 -100
rect -232 -136 -224 -119
rect -207 -136 -199 -119
rect -232 -144 -199 -136
rect -136 -119 -103 -111
rect -79 -113 -64 -100
rect -31 -111 -16 -100
rect -136 -136 -128 -119
rect -111 -136 -103 -119
rect -136 -144 -103 -136
rect -40 -119 -7 -111
rect 16 -113 31 -100
rect 64 -111 79 -100
rect -40 -136 -32 -119
rect -15 -136 -7 -119
rect -40 -144 -7 -136
rect 55 -119 88 -111
rect 112 -113 127 -100
rect 160 -111 175 -100
rect 55 -136 63 -119
rect 80 -136 88 -119
rect 55 -144 88 -136
rect 151 -119 184 -111
rect 208 -113 223 -100
rect 151 -136 159 -119
rect 176 -136 184 -119
rect 151 -144 184 -136
<< polycont >>
rect -176 119 -159 136
rect -80 119 -63 136
rect 15 119 32 136
rect 111 119 128 136
rect 207 119 224 136
rect -224 -136 -207 -119
rect -128 -136 -111 -119
rect -32 -136 -15 -119
rect 63 -136 80 -119
rect 159 -136 176 -119
<< locali >>
rect -305 170 -257 187
rect 257 170 305 187
rect -305 139 -288 170
rect 288 139 305 170
rect -184 119 -176 136
rect -159 119 -151 136
rect -88 119 -80 136
rect -63 119 -55 136
rect 7 119 15 136
rect 32 119 40 136
rect 103 119 111 136
rect 128 119 136 136
rect 199 119 207 136
rect 224 119 232 136
rect -248 94 -231 102
rect -248 -102 -231 -94
rect -200 94 -183 102
rect -200 -102 -183 -94
rect -152 94 -135 102
rect -152 -102 -135 -94
rect -104 94 -87 102
rect -104 -102 -87 -94
rect -56 94 -39 102
rect -56 -102 -39 -94
rect -8 94 9 102
rect -8 -102 9 -94
rect 39 94 56 102
rect 39 -102 56 -94
rect 87 94 104 102
rect 87 -102 104 -94
rect 135 94 152 102
rect 135 -102 152 -94
rect 183 94 200 102
rect 183 -102 200 -94
rect 231 94 248 102
rect 231 -102 248 -94
rect -232 -136 -224 -119
rect -207 -136 -199 -119
rect -136 -136 -128 -119
rect -111 -136 -103 -119
rect -40 -136 -32 -119
rect -15 -136 -7 -119
rect 55 -136 63 -119
rect 80 -136 88 -119
rect 151 -136 159 -119
rect 176 -136 184 -119
rect -305 -170 -288 -139
rect 288 -170 305 -139
rect -305 -187 -257 -170
rect 257 -187 305 -170
<< viali >>
rect -176 119 -159 136
rect -80 119 -63 136
rect 15 119 32 136
rect 111 119 128 136
rect 207 119 224 136
rect -248 -94 -231 94
rect -200 -94 -183 94
rect -152 -94 -135 94
rect -104 -94 -87 94
rect -56 -94 -39 94
rect -8 -94 9 94
rect 39 -94 56 94
rect 87 -94 104 94
rect 135 -94 152 94
rect 183 -94 200 94
rect 231 -94 248 94
rect -224 -136 -207 -119
rect -128 -136 -111 -119
rect -32 -136 -15 -119
rect 63 -136 80 -119
rect 159 -136 176 -119
<< metal1 >>
rect -182 136 -153 139
rect -182 119 -176 136
rect -159 119 -153 136
rect -182 116 -153 119
rect -86 136 -57 139
rect -86 119 -80 136
rect -63 119 -57 136
rect -86 116 -57 119
rect 9 136 38 139
rect 9 119 15 136
rect 32 119 38 136
rect 9 116 38 119
rect 105 136 134 139
rect 105 119 111 136
rect 128 119 134 136
rect 105 116 134 119
rect 201 136 230 139
rect 201 119 207 136
rect 224 119 230 136
rect 201 116 230 119
rect -251 94 -228 100
rect -251 -94 -248 94
rect -231 -94 -228 94
rect -251 -100 -228 -94
rect -203 94 -180 100
rect -203 -94 -200 94
rect -183 -94 -180 94
rect -203 -100 -180 -94
rect -155 94 -132 100
rect -155 -94 -152 94
rect -135 -94 -132 94
rect -155 -100 -132 -94
rect -107 94 -84 100
rect -107 -94 -104 94
rect -87 -94 -84 94
rect -107 -100 -84 -94
rect -59 94 -36 100
rect -59 -94 -56 94
rect -39 -94 -36 94
rect -59 -100 -36 -94
rect -11 94 12 100
rect -11 -94 -8 94
rect 9 -94 12 94
rect -11 -100 12 -94
rect 36 94 59 100
rect 36 -94 39 94
rect 56 -94 59 94
rect 36 -100 59 -94
rect 84 94 107 100
rect 84 -94 87 94
rect 104 -94 107 94
rect 84 -100 107 -94
rect 132 94 155 100
rect 132 -94 135 94
rect 152 -94 155 94
rect 132 -100 155 -94
rect 180 94 203 100
rect 180 -94 183 94
rect 200 -94 203 94
rect 180 -100 203 -94
rect 228 94 251 100
rect 228 -94 231 94
rect 248 -94 251 94
rect 228 -100 251 -94
rect -230 -119 -201 -116
rect -230 -136 -224 -119
rect -207 -136 -201 -119
rect -230 -139 -201 -136
rect -134 -119 -105 -116
rect -134 -136 -128 -119
rect -111 -136 -105 -119
rect -134 -139 -105 -136
rect -38 -119 -9 -116
rect -38 -136 -32 -119
rect -15 -136 -9 -119
rect -38 -139 -9 -136
rect 57 -119 86 -116
rect 57 -136 63 -119
rect 80 -136 86 -119
rect 57 -139 86 -136
rect 153 -119 182 -116
rect 153 -136 159 -119
rect 176 -136 182 -119
rect 153 -139 182 -136
<< properties >>
string FIXED_BBOX -297 -178 297 178
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
