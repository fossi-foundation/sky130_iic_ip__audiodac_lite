magic
tech sky130A
timestamp 1644523392
<< pwell >>
rect -494 -1183 494 1183
<< mvnmos >>
rect -380 54 -330 1054
rect -301 54 -251 1054
rect -222 54 -172 1054
rect -143 54 -93 1054
rect -64 54 -14 1054
rect 15 54 65 1054
rect 94 54 144 1054
rect 173 54 223 1054
rect 252 54 302 1054
rect 331 54 381 1054
rect -380 -1054 -330 -54
rect -301 -1054 -251 -54
rect -222 -1054 -172 -54
rect -143 -1054 -93 -54
rect -64 -1054 -14 -54
rect 15 -1054 65 -54
rect 94 -1054 144 -54
rect 173 -1054 223 -54
rect 252 -1054 302 -54
rect 331 -1054 381 -54
<< mvndiff >>
rect -409 1048 -380 1054
rect -409 60 -403 1048
rect -386 60 -380 1048
rect -409 54 -380 60
rect -330 1048 -301 1054
rect -330 60 -324 1048
rect -307 60 -301 1048
rect -330 54 -301 60
rect -251 1048 -222 1054
rect -251 60 -245 1048
rect -228 60 -222 1048
rect -251 54 -222 60
rect -172 1048 -143 1054
rect -172 60 -166 1048
rect -149 60 -143 1048
rect -172 54 -143 60
rect -93 1048 -64 1054
rect -93 60 -87 1048
rect -70 60 -64 1048
rect -93 54 -64 60
rect -14 1048 15 1054
rect -14 60 -8 1048
rect 9 60 15 1048
rect -14 54 15 60
rect 65 1048 94 1054
rect 65 60 71 1048
rect 88 60 94 1048
rect 65 54 94 60
rect 144 1048 173 1054
rect 144 60 150 1048
rect 167 60 173 1048
rect 144 54 173 60
rect 223 1048 252 1054
rect 223 60 229 1048
rect 246 60 252 1048
rect 223 54 252 60
rect 302 1048 331 1054
rect 302 60 308 1048
rect 325 60 331 1048
rect 302 54 331 60
rect 381 1048 410 1054
rect 381 60 387 1048
rect 404 60 410 1048
rect 381 54 410 60
rect -409 -60 -380 -54
rect -409 -1048 -403 -60
rect -386 -1048 -380 -60
rect -409 -1054 -380 -1048
rect -330 -60 -301 -54
rect -330 -1048 -324 -60
rect -307 -1048 -301 -60
rect -330 -1054 -301 -1048
rect -251 -60 -222 -54
rect -251 -1048 -245 -60
rect -228 -1048 -222 -60
rect -251 -1054 -222 -1048
rect -172 -60 -143 -54
rect -172 -1048 -166 -60
rect -149 -1048 -143 -60
rect -172 -1054 -143 -1048
rect -93 -60 -64 -54
rect -93 -1048 -87 -60
rect -70 -1048 -64 -60
rect -93 -1054 -64 -1048
rect -14 -60 15 -54
rect -14 -1048 -8 -60
rect 9 -1048 15 -60
rect -14 -1054 15 -1048
rect 65 -60 94 -54
rect 65 -1048 71 -60
rect 88 -1048 94 -60
rect 65 -1054 94 -1048
rect 144 -60 173 -54
rect 144 -1048 150 -60
rect 167 -1048 173 -60
rect 144 -1054 173 -1048
rect 223 -60 252 -54
rect 223 -1048 229 -60
rect 246 -1048 252 -60
rect 223 -1054 252 -1048
rect 302 -60 331 -54
rect 302 -1048 308 -60
rect 325 -1048 331 -60
rect 302 -1054 331 -1048
rect 381 -60 410 -54
rect 381 -1048 387 -60
rect 404 -1048 410 -60
rect 381 -1054 410 -1048
<< mvndiffc >>
rect -403 60 -386 1048
rect -324 60 -307 1048
rect -245 60 -228 1048
rect -166 60 -149 1048
rect -87 60 -70 1048
rect -8 60 9 1048
rect 71 60 88 1048
rect 150 60 167 1048
rect 229 60 246 1048
rect 308 60 325 1048
rect 387 60 404 1048
rect -403 -1048 -386 -60
rect -324 -1048 -307 -60
rect -245 -1048 -228 -60
rect -166 -1048 -149 -60
rect -87 -1048 -70 -60
rect -8 -1048 9 -60
rect 71 -1048 88 -60
rect 150 -1048 167 -60
rect 229 -1048 246 -60
rect 308 -1048 325 -60
rect 387 -1048 404 -60
<< mvpsubdiff >>
rect -476 1159 476 1165
rect -476 1142 -422 1159
rect 422 1142 476 1159
rect -476 1136 476 1142
rect -476 1111 -447 1136
rect -476 -1111 -470 1111
rect -453 -1111 -447 1111
rect 447 1111 476 1136
rect -476 -1136 -447 -1111
rect 447 -1111 453 1111
rect 470 -1111 476 1111
rect 447 -1136 476 -1111
rect -476 -1142 476 -1136
rect -476 -1159 -422 -1142
rect 422 -1159 476 -1142
rect -476 -1165 476 -1159
<< mvpsubdiffcont >>
rect -422 1142 422 1159
rect -470 -1111 -453 1111
rect 453 -1111 470 1111
rect -422 -1159 422 -1142
<< poly >>
rect -380 1090 -330 1098
rect -380 1073 -372 1090
rect -338 1073 -330 1090
rect -380 1054 -330 1073
rect -301 1090 -251 1098
rect -301 1073 -293 1090
rect -259 1073 -251 1090
rect -301 1054 -251 1073
rect -222 1090 -172 1098
rect -222 1073 -214 1090
rect -180 1073 -172 1090
rect -222 1054 -172 1073
rect -143 1090 -93 1098
rect -143 1073 -135 1090
rect -101 1073 -93 1090
rect -143 1054 -93 1073
rect -64 1090 -14 1098
rect -64 1073 -56 1090
rect -22 1073 -14 1090
rect -64 1054 -14 1073
rect 15 1090 65 1098
rect 15 1073 23 1090
rect 57 1073 65 1090
rect 15 1054 65 1073
rect 94 1090 144 1098
rect 94 1073 102 1090
rect 136 1073 144 1090
rect 94 1054 144 1073
rect 173 1090 223 1098
rect 173 1073 181 1090
rect 215 1073 223 1090
rect 173 1054 223 1073
rect 252 1090 302 1098
rect 252 1073 260 1090
rect 294 1073 302 1090
rect 252 1054 302 1073
rect 331 1090 381 1098
rect 331 1073 339 1090
rect 373 1073 381 1090
rect 331 1054 381 1073
rect -380 35 -330 54
rect -380 18 -372 35
rect -338 18 -330 35
rect -380 -18 -330 18
rect -380 -35 -372 -18
rect -338 -35 -330 -18
rect -380 -54 -330 -35
rect -301 35 -251 54
rect -301 18 -293 35
rect -259 18 -251 35
rect -301 -18 -251 18
rect -301 -35 -293 -18
rect -259 -35 -251 -18
rect -301 -54 -251 -35
rect -222 35 -172 54
rect -222 18 -214 35
rect -180 18 -172 35
rect -222 -18 -172 18
rect -222 -35 -214 -18
rect -180 -35 -172 -18
rect -222 -54 -172 -35
rect -143 35 -93 54
rect -143 18 -135 35
rect -101 18 -93 35
rect -143 -18 -93 18
rect -143 -35 -135 -18
rect -101 -35 -93 -18
rect -143 -54 -93 -35
rect -64 35 -14 54
rect -64 18 -56 35
rect -22 18 -14 35
rect -64 -18 -14 18
rect -64 -35 -56 -18
rect -22 -35 -14 -18
rect -64 -54 -14 -35
rect 15 35 65 54
rect 15 18 23 35
rect 57 18 65 35
rect 15 -18 65 18
rect 15 -35 23 -18
rect 57 -35 65 -18
rect 15 -54 65 -35
rect 94 35 144 54
rect 94 18 102 35
rect 136 18 144 35
rect 94 -18 144 18
rect 94 -35 102 -18
rect 136 -35 144 -18
rect 94 -54 144 -35
rect 173 35 223 54
rect 173 18 181 35
rect 215 18 223 35
rect 173 -18 223 18
rect 173 -35 181 -18
rect 215 -35 223 -18
rect 173 -54 223 -35
rect 252 35 302 54
rect 252 18 260 35
rect 294 18 302 35
rect 252 -18 302 18
rect 252 -35 260 -18
rect 294 -35 302 -18
rect 252 -54 302 -35
rect 331 35 381 54
rect 331 18 339 35
rect 373 18 381 35
rect 331 -18 381 18
rect 331 -35 339 -18
rect 373 -35 381 -18
rect 331 -54 381 -35
rect -380 -1073 -330 -1054
rect -380 -1090 -372 -1073
rect -338 -1090 -330 -1073
rect -380 -1098 -330 -1090
rect -301 -1073 -251 -1054
rect -301 -1090 -293 -1073
rect -259 -1090 -251 -1073
rect -301 -1098 -251 -1090
rect -222 -1073 -172 -1054
rect -222 -1090 -214 -1073
rect -180 -1090 -172 -1073
rect -222 -1098 -172 -1090
rect -143 -1073 -93 -1054
rect -143 -1090 -135 -1073
rect -101 -1090 -93 -1073
rect -143 -1098 -93 -1090
rect -64 -1073 -14 -1054
rect -64 -1090 -56 -1073
rect -22 -1090 -14 -1073
rect -64 -1098 -14 -1090
rect 15 -1073 65 -1054
rect 15 -1090 23 -1073
rect 57 -1090 65 -1073
rect 15 -1098 65 -1090
rect 94 -1073 144 -1054
rect 94 -1090 102 -1073
rect 136 -1090 144 -1073
rect 94 -1098 144 -1090
rect 173 -1073 223 -1054
rect 173 -1090 181 -1073
rect 215 -1090 223 -1073
rect 173 -1098 223 -1090
rect 252 -1073 302 -1054
rect 252 -1090 260 -1073
rect 294 -1090 302 -1073
rect 252 -1098 302 -1090
rect 331 -1073 381 -1054
rect 331 -1090 339 -1073
rect 373 -1090 381 -1073
rect 331 -1098 381 -1090
<< polycont >>
rect -372 1073 -338 1090
rect -293 1073 -259 1090
rect -214 1073 -180 1090
rect -135 1073 -101 1090
rect -56 1073 -22 1090
rect 23 1073 57 1090
rect 102 1073 136 1090
rect 181 1073 215 1090
rect 260 1073 294 1090
rect 339 1073 373 1090
rect -372 18 -338 35
rect -372 -35 -338 -18
rect -293 18 -259 35
rect -293 -35 -259 -18
rect -214 18 -180 35
rect -214 -35 -180 -18
rect -135 18 -101 35
rect -135 -35 -101 -18
rect -56 18 -22 35
rect -56 -35 -22 -18
rect 23 18 57 35
rect 23 -35 57 -18
rect 102 18 136 35
rect 102 -35 136 -18
rect 181 18 215 35
rect 181 -35 215 -18
rect 260 18 294 35
rect 260 -35 294 -18
rect 339 18 373 35
rect 339 -35 373 -18
rect -372 -1090 -338 -1073
rect -293 -1090 -259 -1073
rect -214 -1090 -180 -1073
rect -135 -1090 -101 -1073
rect -56 -1090 -22 -1073
rect 23 -1090 57 -1073
rect 102 -1090 136 -1073
rect 181 -1090 215 -1073
rect 260 -1090 294 -1073
rect 339 -1090 373 -1073
<< locali >>
rect -470 1142 -422 1159
rect 422 1142 470 1159
rect -470 1111 -453 1142
rect 453 1111 470 1142
rect -380 1073 -372 1090
rect -338 1073 -330 1090
rect -301 1073 -293 1090
rect -259 1073 -251 1090
rect -222 1073 -214 1090
rect -180 1073 -172 1090
rect -143 1073 -135 1090
rect -101 1073 -93 1090
rect -64 1073 -56 1090
rect -22 1073 -14 1090
rect 15 1073 23 1090
rect 57 1073 65 1090
rect 94 1073 102 1090
rect 136 1073 144 1090
rect 173 1073 181 1090
rect 215 1073 223 1090
rect 252 1073 260 1090
rect 294 1073 302 1090
rect 331 1073 339 1090
rect 373 1073 381 1090
rect -403 1048 -386 1056
rect -403 52 -386 60
rect -324 1048 -307 1056
rect -324 52 -307 60
rect -245 1048 -228 1056
rect -245 52 -228 60
rect -166 1048 -149 1056
rect -166 52 -149 60
rect -87 1048 -70 1056
rect -87 52 -70 60
rect -8 1048 9 1056
rect -8 52 9 60
rect 71 1048 88 1056
rect 71 52 88 60
rect 150 1048 167 1056
rect 150 52 167 60
rect 229 1048 246 1056
rect 229 52 246 60
rect 308 1048 325 1056
rect 308 52 325 60
rect 387 1048 404 1056
rect 387 52 404 60
rect -380 18 -372 35
rect -338 18 -330 35
rect -301 18 -293 35
rect -259 18 -251 35
rect -222 18 -214 35
rect -180 18 -172 35
rect -143 18 -135 35
rect -101 18 -93 35
rect -64 18 -56 35
rect -22 18 -14 35
rect 15 18 23 35
rect 57 18 65 35
rect 94 18 102 35
rect 136 18 144 35
rect 173 18 181 35
rect 215 18 223 35
rect 252 18 260 35
rect 294 18 302 35
rect 331 18 339 35
rect 373 18 381 35
rect -380 -35 -372 -18
rect -338 -35 -330 -18
rect -301 -35 -293 -18
rect -259 -35 -251 -18
rect -222 -35 -214 -18
rect -180 -35 -172 -18
rect -143 -35 -135 -18
rect -101 -35 -93 -18
rect -64 -35 -56 -18
rect -22 -35 -14 -18
rect 15 -35 23 -18
rect 57 -35 65 -18
rect 94 -35 102 -18
rect 136 -35 144 -18
rect 173 -35 181 -18
rect 215 -35 223 -18
rect 252 -35 260 -18
rect 294 -35 302 -18
rect 331 -35 339 -18
rect 373 -35 381 -18
rect -403 -60 -386 -52
rect -403 -1056 -386 -1048
rect -324 -60 -307 -52
rect -324 -1056 -307 -1048
rect -245 -60 -228 -52
rect -245 -1056 -228 -1048
rect -166 -60 -149 -52
rect -166 -1056 -149 -1048
rect -87 -60 -70 -52
rect -87 -1056 -70 -1048
rect -8 -60 9 -52
rect -8 -1056 9 -1048
rect 71 -60 88 -52
rect 71 -1056 88 -1048
rect 150 -60 167 -52
rect 150 -1056 167 -1048
rect 229 -60 246 -52
rect 229 -1056 246 -1048
rect 308 -60 325 -52
rect 308 -1056 325 -1048
rect 387 -60 404 -52
rect 387 -1056 404 -1048
rect -380 -1090 -372 -1073
rect -338 -1090 -330 -1073
rect -301 -1090 -293 -1073
rect -259 -1090 -251 -1073
rect -222 -1090 -214 -1073
rect -180 -1090 -172 -1073
rect -143 -1090 -135 -1073
rect -101 -1090 -93 -1073
rect -64 -1090 -56 -1073
rect -22 -1090 -14 -1073
rect 15 -1090 23 -1073
rect 57 -1090 65 -1073
rect 94 -1090 102 -1073
rect 136 -1090 144 -1073
rect 173 -1090 181 -1073
rect 215 -1090 223 -1073
rect 252 -1090 260 -1073
rect 294 -1090 302 -1073
rect 331 -1090 339 -1073
rect 373 -1090 381 -1073
rect -470 -1142 -453 -1111
rect 453 -1142 470 -1111
rect -470 -1159 -422 -1142
rect 422 -1159 470 -1142
<< viali >>
rect -372 1073 -338 1090
rect -293 1073 -259 1090
rect -214 1073 -180 1090
rect -135 1073 -101 1090
rect -56 1073 -22 1090
rect 23 1073 57 1090
rect 102 1073 136 1090
rect 181 1073 215 1090
rect 260 1073 294 1090
rect 339 1073 373 1090
rect -403 60 -386 1048
rect -324 60 -307 1048
rect -245 60 -228 1048
rect -166 60 -149 1048
rect -87 60 -70 1048
rect -8 60 9 1048
rect 71 60 88 1048
rect 150 60 167 1048
rect 229 60 246 1048
rect 308 60 325 1048
rect 387 60 404 1048
rect -372 18 -338 35
rect -293 18 -259 35
rect -214 18 -180 35
rect -135 18 -101 35
rect -56 18 -22 35
rect 23 18 57 35
rect 102 18 136 35
rect 181 18 215 35
rect 260 18 294 35
rect 339 18 373 35
rect -372 -35 -338 -18
rect -293 -35 -259 -18
rect -214 -35 -180 -18
rect -135 -35 -101 -18
rect -56 -35 -22 -18
rect 23 -35 57 -18
rect 102 -35 136 -18
rect 181 -35 215 -18
rect 260 -35 294 -18
rect 339 -35 373 -18
rect -403 -1048 -386 -60
rect -324 -1048 -307 -60
rect -245 -1048 -228 -60
rect -166 -1048 -149 -60
rect -87 -1048 -70 -60
rect -8 -1048 9 -60
rect 71 -1048 88 -60
rect 150 -1048 167 -60
rect 229 -1048 246 -60
rect 308 -1048 325 -60
rect 387 -1048 404 -60
rect -372 -1090 -338 -1073
rect -293 -1090 -259 -1073
rect -214 -1090 -180 -1073
rect -135 -1090 -101 -1073
rect -56 -1090 -22 -1073
rect 23 -1090 57 -1073
rect 102 -1090 136 -1073
rect 181 -1090 215 -1073
rect 260 -1090 294 -1073
rect 339 -1090 373 -1073
<< metal1 >>
rect -378 1090 -332 1093
rect -378 1073 -372 1090
rect -338 1073 -332 1090
rect -378 1070 -332 1073
rect -299 1090 -253 1093
rect -299 1073 -293 1090
rect -259 1073 -253 1090
rect -299 1070 -253 1073
rect -220 1090 -174 1093
rect -220 1073 -214 1090
rect -180 1073 -174 1090
rect -220 1070 -174 1073
rect -141 1090 -95 1093
rect -141 1073 -135 1090
rect -101 1073 -95 1090
rect -141 1070 -95 1073
rect -62 1090 -16 1093
rect -62 1073 -56 1090
rect -22 1073 -16 1090
rect -62 1070 -16 1073
rect 17 1090 63 1093
rect 17 1073 23 1090
rect 57 1073 63 1090
rect 17 1070 63 1073
rect 96 1090 142 1093
rect 96 1073 102 1090
rect 136 1073 142 1090
rect 96 1070 142 1073
rect 175 1090 221 1093
rect 175 1073 181 1090
rect 215 1073 221 1090
rect 175 1070 221 1073
rect 254 1090 300 1093
rect 254 1073 260 1090
rect 294 1073 300 1090
rect 254 1070 300 1073
rect 333 1090 379 1093
rect 333 1073 339 1090
rect 373 1073 379 1090
rect 333 1070 379 1073
rect -406 1048 -383 1054
rect -406 60 -403 1048
rect -386 60 -383 1048
rect -406 54 -383 60
rect -327 1048 -304 1054
rect -327 60 -324 1048
rect -307 60 -304 1048
rect -327 54 -304 60
rect -248 1048 -225 1054
rect -248 60 -245 1048
rect -228 60 -225 1048
rect -248 54 -225 60
rect -169 1048 -146 1054
rect -169 60 -166 1048
rect -149 60 -146 1048
rect -169 54 -146 60
rect -90 1048 -67 1054
rect -90 60 -87 1048
rect -70 60 -67 1048
rect -90 54 -67 60
rect -11 1048 12 1054
rect -11 60 -8 1048
rect 9 60 12 1048
rect -11 54 12 60
rect 68 1048 91 1054
rect 68 60 71 1048
rect 88 60 91 1048
rect 68 54 91 60
rect 147 1048 170 1054
rect 147 60 150 1048
rect 167 60 170 1048
rect 147 54 170 60
rect 226 1048 249 1054
rect 226 60 229 1048
rect 246 60 249 1048
rect 226 54 249 60
rect 305 1048 328 1054
rect 305 60 308 1048
rect 325 60 328 1048
rect 305 54 328 60
rect 384 1048 407 1054
rect 384 60 387 1048
rect 404 60 407 1048
rect 384 54 407 60
rect -378 35 -332 38
rect -378 18 -372 35
rect -338 18 -332 35
rect -378 15 -332 18
rect -299 35 -253 38
rect -299 18 -293 35
rect -259 18 -253 35
rect -299 15 -253 18
rect -220 35 -174 38
rect -220 18 -214 35
rect -180 18 -174 35
rect -220 15 -174 18
rect -141 35 -95 38
rect -141 18 -135 35
rect -101 18 -95 35
rect -141 15 -95 18
rect -62 35 -16 38
rect -62 18 -56 35
rect -22 18 -16 35
rect -62 15 -16 18
rect 17 35 63 38
rect 17 18 23 35
rect 57 18 63 35
rect 17 15 63 18
rect 96 35 142 38
rect 96 18 102 35
rect 136 18 142 35
rect 96 15 142 18
rect 175 35 221 38
rect 175 18 181 35
rect 215 18 221 35
rect 175 15 221 18
rect 254 35 300 38
rect 254 18 260 35
rect 294 18 300 35
rect 254 15 300 18
rect 333 35 379 38
rect 333 18 339 35
rect 373 18 379 35
rect 333 15 379 18
rect -378 -18 -332 -15
rect -378 -35 -372 -18
rect -338 -35 -332 -18
rect -378 -38 -332 -35
rect -299 -18 -253 -15
rect -299 -35 -293 -18
rect -259 -35 -253 -18
rect -299 -38 -253 -35
rect -220 -18 -174 -15
rect -220 -35 -214 -18
rect -180 -35 -174 -18
rect -220 -38 -174 -35
rect -141 -18 -95 -15
rect -141 -35 -135 -18
rect -101 -35 -95 -18
rect -141 -38 -95 -35
rect -62 -18 -16 -15
rect -62 -35 -56 -18
rect -22 -35 -16 -18
rect -62 -38 -16 -35
rect 17 -18 63 -15
rect 17 -35 23 -18
rect 57 -35 63 -18
rect 17 -38 63 -35
rect 96 -18 142 -15
rect 96 -35 102 -18
rect 136 -35 142 -18
rect 96 -38 142 -35
rect 175 -18 221 -15
rect 175 -35 181 -18
rect 215 -35 221 -18
rect 175 -38 221 -35
rect 254 -18 300 -15
rect 254 -35 260 -18
rect 294 -35 300 -18
rect 254 -38 300 -35
rect 333 -18 379 -15
rect 333 -35 339 -18
rect 373 -35 379 -18
rect 333 -38 379 -35
rect -406 -60 -383 -54
rect -406 -1048 -403 -60
rect -386 -1048 -383 -60
rect -406 -1054 -383 -1048
rect -327 -60 -304 -54
rect -327 -1048 -324 -60
rect -307 -1048 -304 -60
rect -327 -1054 -304 -1048
rect -248 -60 -225 -54
rect -248 -1048 -245 -60
rect -228 -1048 -225 -60
rect -248 -1054 -225 -1048
rect -169 -60 -146 -54
rect -169 -1048 -166 -60
rect -149 -1048 -146 -60
rect -169 -1054 -146 -1048
rect -90 -60 -67 -54
rect -90 -1048 -87 -60
rect -70 -1048 -67 -60
rect -90 -1054 -67 -1048
rect -11 -60 12 -54
rect -11 -1048 -8 -60
rect 9 -1048 12 -60
rect -11 -1054 12 -1048
rect 68 -60 91 -54
rect 68 -1048 71 -60
rect 88 -1048 91 -60
rect 68 -1054 91 -1048
rect 147 -60 170 -54
rect 147 -1048 150 -60
rect 167 -1048 170 -60
rect 147 -1054 170 -1048
rect 226 -60 249 -54
rect 226 -1048 229 -60
rect 246 -1048 249 -60
rect 226 -1054 249 -1048
rect 305 -60 328 -54
rect 305 -1048 308 -60
rect 325 -1048 328 -60
rect 305 -1054 328 -1048
rect 384 -60 407 -54
rect 384 -1048 387 -60
rect 404 -1048 407 -60
rect 384 -1054 407 -1048
rect -378 -1073 -332 -1070
rect -378 -1090 -372 -1073
rect -338 -1090 -332 -1073
rect -378 -1093 -332 -1090
rect -299 -1073 -253 -1070
rect -299 -1090 -293 -1073
rect -259 -1090 -253 -1073
rect -299 -1093 -253 -1090
rect -220 -1073 -174 -1070
rect -220 -1090 -214 -1073
rect -180 -1090 -174 -1073
rect -220 -1093 -174 -1090
rect -141 -1073 -95 -1070
rect -141 -1090 -135 -1073
rect -101 -1090 -95 -1073
rect -141 -1093 -95 -1090
rect -62 -1073 -16 -1070
rect -62 -1090 -56 -1073
rect -22 -1090 -16 -1073
rect -62 -1093 -16 -1090
rect 17 -1073 63 -1070
rect 17 -1090 23 -1073
rect 57 -1090 63 -1073
rect 17 -1093 63 -1090
rect 96 -1073 142 -1070
rect 96 -1090 102 -1073
rect 136 -1090 142 -1073
rect 96 -1093 142 -1090
rect 175 -1073 221 -1070
rect 175 -1090 181 -1073
rect 215 -1090 221 -1073
rect 175 -1093 221 -1090
rect 254 -1073 300 -1070
rect 254 -1090 260 -1073
rect 294 -1090 300 -1073
rect 254 -1093 300 -1090
rect 333 -1073 379 -1070
rect 333 -1090 339 -1073
rect 373 -1090 379 -1073
rect 333 -1093 379 -1090
<< properties >>
string FIXED_BBOX -462 -1151 462 1151
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 0.5 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
