magic
tech sky130A
timestamp 1721163516
<< pwell >>
rect -297 -629 297 629
<< mvnmos >>
rect -183 -500 -133 500
rect -104 -500 -54 500
rect -25 -500 25 500
rect 54 -500 104 500
rect 133 -500 183 500
<< mvndiff >>
rect -212 494 -183 500
rect -212 -494 -206 494
rect -189 -494 -183 494
rect -212 -500 -183 -494
rect -133 494 -104 500
rect -133 -494 -127 494
rect -110 -494 -104 494
rect -133 -500 -104 -494
rect -54 494 -25 500
rect -54 -494 -48 494
rect -31 -494 -25 494
rect -54 -500 -25 -494
rect 25 494 54 500
rect 25 -494 31 494
rect 48 -494 54 494
rect 25 -500 54 -494
rect 104 494 133 500
rect 104 -494 110 494
rect 127 -494 133 494
rect 104 -500 133 -494
rect 183 494 212 500
rect 183 -494 189 494
rect 206 -494 212 494
rect 183 -500 212 -494
<< mvndiffc >>
rect -206 -494 -189 494
rect -127 -494 -110 494
rect -48 -494 -31 494
rect 31 -494 48 494
rect 110 -494 127 494
rect 189 -494 206 494
<< mvpsubdiff >>
rect -279 605 279 611
rect -279 588 -225 605
rect 225 588 279 605
rect -279 582 279 588
rect -279 557 -250 582
rect -279 -557 -273 557
rect -256 -557 -250 557
rect 250 557 279 582
rect -279 -582 -250 -557
rect 250 -557 256 557
rect 273 -557 279 557
rect 250 -582 279 -557
rect -279 -588 279 -582
rect -279 -605 -225 -588
rect 225 -605 279 -588
rect -279 -611 279 -605
<< mvpsubdiffcont >>
rect -225 588 225 605
rect -273 -557 -256 557
rect 256 -557 273 557
rect -225 -605 225 -588
<< poly >>
rect -183 536 -133 544
rect -183 519 -175 536
rect -141 519 -133 536
rect -183 500 -133 519
rect -104 536 -54 544
rect -104 519 -96 536
rect -62 519 -54 536
rect -104 500 -54 519
rect -25 536 25 544
rect -25 519 -17 536
rect 17 519 25 536
rect -25 500 25 519
rect 54 536 104 544
rect 54 519 62 536
rect 96 519 104 536
rect 54 500 104 519
rect 133 536 183 544
rect 133 519 141 536
rect 175 519 183 536
rect 133 500 183 519
rect -183 -519 -133 -500
rect -183 -536 -175 -519
rect -141 -536 -133 -519
rect -183 -544 -133 -536
rect -104 -519 -54 -500
rect -104 -536 -96 -519
rect -62 -536 -54 -519
rect -104 -544 -54 -536
rect -25 -519 25 -500
rect -25 -536 -17 -519
rect 17 -536 25 -519
rect -25 -544 25 -536
rect 54 -519 104 -500
rect 54 -536 62 -519
rect 96 -536 104 -519
rect 54 -544 104 -536
rect 133 -519 183 -500
rect 133 -536 141 -519
rect 175 -536 183 -519
rect 133 -544 183 -536
<< polycont >>
rect -175 519 -141 536
rect -96 519 -62 536
rect -17 519 17 536
rect 62 519 96 536
rect 141 519 175 536
rect -175 -536 -141 -519
rect -96 -536 -62 -519
rect -17 -536 17 -519
rect 62 -536 96 -519
rect 141 -536 175 -519
<< locali >>
rect -273 588 -225 605
rect 225 588 273 605
rect -273 557 -256 588
rect 256 557 273 588
rect -183 519 -175 536
rect -141 519 -133 536
rect -104 519 -96 536
rect -62 519 -54 536
rect -25 519 -17 536
rect 17 519 25 536
rect 54 519 62 536
rect 96 519 104 536
rect 133 519 141 536
rect 175 519 183 536
rect -206 494 -189 502
rect -206 -502 -189 -494
rect -127 494 -110 502
rect -127 -502 -110 -494
rect -48 494 -31 502
rect -48 -502 -31 -494
rect 31 494 48 502
rect 31 -502 48 -494
rect 110 494 127 502
rect 110 -502 127 -494
rect 189 494 206 502
rect 189 -502 206 -494
rect -183 -536 -175 -519
rect -141 -536 -133 -519
rect -104 -536 -96 -519
rect -62 -536 -54 -519
rect -25 -536 -17 -519
rect 17 -536 25 -519
rect 54 -536 62 -519
rect 96 -536 104 -519
rect 133 -536 141 -519
rect 175 -536 183 -519
rect -273 -588 -256 -557
rect 256 -588 273 -557
rect -273 -605 -225 -588
rect 225 -605 273 -588
<< viali >>
rect -175 519 -141 536
rect -96 519 -62 536
rect -17 519 17 536
rect 62 519 96 536
rect 141 519 175 536
rect -206 -494 -189 494
rect -127 -494 -110 494
rect -48 -494 -31 494
rect 31 -494 48 494
rect 110 -494 127 494
rect 189 -494 206 494
rect -175 -536 -141 -519
rect -96 -536 -62 -519
rect -17 -536 17 -519
rect 62 -536 96 -519
rect 141 -536 175 -519
<< metal1 >>
rect -181 536 -135 539
rect -181 519 -175 536
rect -141 519 -135 536
rect -181 516 -135 519
rect -102 536 -56 539
rect -102 519 -96 536
rect -62 519 -56 536
rect -102 516 -56 519
rect -23 536 23 539
rect -23 519 -17 536
rect 17 519 23 536
rect -23 516 23 519
rect 56 536 102 539
rect 56 519 62 536
rect 96 519 102 536
rect 56 516 102 519
rect 135 536 181 539
rect 135 519 141 536
rect 175 519 181 536
rect 135 516 181 519
rect -209 494 -186 500
rect -209 -494 -206 494
rect -189 -494 -186 494
rect -209 -500 -186 -494
rect -130 494 -107 500
rect -130 -494 -127 494
rect -110 -494 -107 494
rect -130 -500 -107 -494
rect -51 494 -28 500
rect -51 -494 -48 494
rect -31 -494 -28 494
rect -51 -500 -28 -494
rect 28 494 51 500
rect 28 -494 31 494
rect 48 -494 51 494
rect 28 -500 51 -494
rect 107 494 130 500
rect 107 -494 110 494
rect 127 -494 130 494
rect 107 -500 130 -494
rect 186 494 209 500
rect 186 -494 189 494
rect 206 -494 209 494
rect 186 -500 209 -494
rect -181 -519 -135 -516
rect -181 -536 -175 -519
rect -141 -536 -135 -519
rect -181 -539 -135 -536
rect -102 -519 -56 -516
rect -102 -536 -96 -519
rect -62 -536 -56 -519
rect -102 -539 -56 -536
rect -23 -519 23 -516
rect -23 -536 -17 -519
rect 17 -536 23 -519
rect -23 -539 23 -536
rect 56 -519 102 -516
rect 56 -536 62 -519
rect 96 -536 102 -519
rect 56 -539 102 -536
rect 135 -519 181 -516
rect 135 -536 141 -519
rect 175 -536 181 -519
rect 135 -539 181 -536
<< properties >>
string FIXED_BBOX -264 -596 264 596
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.50 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
