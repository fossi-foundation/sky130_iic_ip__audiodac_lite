magic
tech sky130A
magscale 1 2
timestamp 1747753680
<< dnwell >>
rect -206 -190 14946 28568
<< nwell >>
rect -316 28362 15056 28678
rect -316 16792 47 28362
rect 2533 28114 2853 28362
rect 2521 28094 2853 28114
rect 2521 27358 2811 28094
rect 2541 26124 2809 27358
rect 2541 24140 2807 26124
rect 2527 23558 2849 24140
rect 2527 23536 3061 23558
rect 2551 23530 3061 23536
rect 14720 19064 15056 28362
rect -316 11594 0 16792
rect -316 16 27 11594
rect 14740 9302 15056 19064
rect 2529 4836 2621 4838
rect 2529 4818 3047 4836
rect 2529 4808 2833 4818
rect 2495 1242 2833 4808
rect 2501 218 2833 1242
rect 2501 46 2897 218
rect 2435 16 2969 46
rect 14720 16 15056 9302
rect -316 -300 15056 16
<< mvnsubdiff >>
rect -249 28591 14989 28611
rect -249 28557 -169 28591
rect 14909 28557 14989 28591
rect -249 28537 14989 28557
rect -249 28531 -175 28537
rect -249 -153 -229 28531
rect -195 -153 -175 28531
rect -249 -159 -175 -153
rect 14915 28531 14989 28537
rect 14915 -153 14935 28531
rect 14969 -153 14989 28531
rect 14915 -159 14989 -153
rect -249 -179 14989 -159
rect -249 -213 -169 -179
rect 14909 -213 14989 -179
rect -249 -233 14989 -213
<< mvnsubdiffcont >>
rect -169 28557 14909 28591
rect -229 -153 -195 28531
rect 14935 -153 14969 28531
rect -169 -213 14909 -179
<< locali >>
rect -249 28591 14991 28621
rect -249 28557 -169 28591
rect 14909 28557 14991 28591
rect -249 28531 14991 28557
rect -249 -153 -229 28531
rect -195 28503 14935 28531
rect -195 -139 -131 28503
rect 117 10632 257 11300
rect 2297 11280 2445 11302
rect 121 304 255 10632
rect 2297 342 2449 11280
rect 121 298 273 304
rect 123 292 273 298
rect 2297 292 2451 342
rect 14873 -139 14935 28503
rect -195 -153 14935 -139
rect 14969 -153 14991 28531
rect -249 -179 14991 -153
rect -249 -213 -169 -179
rect 14909 -213 14991 -179
rect -249 -257 14991 -213
<< metal1 >>
rect -249 28503 14991 28621
rect -249 25235 -131 28503
rect -249 25232 276 25235
rect -249 23206 267 25232
rect 2341 23206 2351 25232
rect -249 23202 276 23206
rect -249 5650 -131 23202
rect 3343 21278 3349 21386
rect 3457 21278 3463 21386
rect 2738 18784 2965 18974
rect 293 16928 303 17048
rect 2301 16928 2311 17048
rect 2738 15727 2928 18784
rect 2738 15537 3386 15727
rect 1 12929 103 15196
rect 3196 13773 3386 15537
rect 3196 13583 3660 13773
rect 4349 13604 4787 13764
rect 4627 12132 4787 13604
rect 3929 11972 4787 12132
rect 3929 11956 4089 11972
rect 2775 11796 4089 11956
rect 275 11346 285 11440
rect 2285 11346 2295 11440
rect 2775 9236 2935 11796
rect 3343 6934 3349 7042
rect 3457 6934 3463 7042
rect 229 5650 239 5652
rect -249 3682 239 5650
rect -249 -139 -131 3682
rect 229 3680 239 3682
rect 2335 3680 2345 5652
rect 14873 -139 14991 28503
rect -249 -257 14991 -139
<< via1 >>
rect 267 23206 2341 25232
rect 3349 21278 3457 21386
rect 303 16928 2301 17048
rect 285 11346 2285 11440
rect 3349 6934 3457 7042
rect 239 3680 2335 5652
<< metal2 >>
rect 267 25232 2341 25242
rect 267 23196 2341 23206
rect 3349 21386 3457 21392
rect 3340 21278 3349 21386
rect 3457 21278 3466 21386
rect 3349 21272 3457 21278
rect 4979 19890 5079 19899
rect 4979 19721 5079 19730
rect 299 17048 5021 17468
rect 299 16928 303 17048
rect 2301 16928 5021 17048
rect 299 16852 5021 16928
rect 2546 16057 2610 16091
rect 2546 16056 2721 16057
rect 2546 15975 2831 16056
rect 2546 15971 2610 15975
rect 2721 15917 2831 15975
rect 4574 15960 4744 15969
rect 3886 15917 3968 15960
rect 2721 15836 3968 15917
rect 2831 15835 3968 15836
rect 973 15701 982 15799
rect 1080 15701 1089 15799
rect 2124 15789 2222 15798
rect 3886 15790 3968 15835
rect 4200 15790 4574 15960
rect 4574 15781 4744 15790
rect 2124 15682 2222 15691
rect 3570 12536 3834 12576
rect 3095 12412 4987 12536
rect 3095 12286 3219 12412
rect 3570 12406 3834 12412
rect 544 12161 684 12285
rect 2665 12162 3219 12286
rect 4863 11540 4987 12412
rect 277 11440 5045 11540
rect 277 11346 285 11440
rect 2285 11346 5045 11440
rect 277 11152 5045 11346
rect 3349 7042 3457 7048
rect 3340 6934 3349 7042
rect 3457 6934 3466 7042
rect 3349 6928 3457 6934
rect 239 5652 2335 5662
rect 239 3670 2335 3680
<< via2 >>
rect 267 23206 2341 25232
rect 3349 21278 3457 21386
rect 982 15701 1080 15799
rect 4574 15790 4744 15960
rect 2124 15691 2222 15789
rect 3349 6934 3457 7042
rect 239 3680 2335 5652
<< metal3 >>
rect 267 25237 8465 25260
rect 257 25232 8465 25237
rect 257 23206 267 25232
rect 2341 23206 8465 25232
rect 257 23201 2351 23206
rect 8699 21846 12023 26696
rect 3344 21386 3462 21391
rect 2809 21278 3349 21386
rect 3457 21278 3462 21386
rect 2809 16150 2917 21278
rect 3344 21273 3462 21278
rect 8699 21046 12031 21846
rect 12481 21092 14317 22848
rect 977 16042 2917 16150
rect 5433 19650 8517 19712
rect 977 15799 1085 16042
rect 5433 15966 5477 19650
rect 977 15701 982 15799
rect 1080 15701 1085 15799
rect 4563 15960 5477 15966
rect 977 15688 1085 15701
rect 2119 15789 3165 15794
rect 2119 15691 2124 15789
rect 2222 15691 3165 15789
rect 4563 15790 4574 15960
rect 4744 15790 5477 15960
rect 4563 15780 5477 15790
rect 2119 15686 3165 15691
rect 70 12509 2750 12589
rect 70 12329 360 12409
rect 3057 12006 3165 15686
rect 2811 11898 3165 12006
rect 5433 15100 5477 15780
rect 8439 15100 8517 19650
rect 8707 16610 12031 21046
rect 2811 7042 2919 11898
rect 3344 7042 3462 7047
rect 2811 6934 3349 7042
rect 3457 6934 3462 7042
rect 3344 6929 3462 6934
rect 5433 6526 8517 15100
rect 8703 16196 12031 16610
rect 8703 13336 12027 16196
rect 8703 11358 8833 13336
rect 229 5652 8449 5662
rect 229 3680 239 5652
rect 2335 3680 8449 5652
rect 229 3676 8449 3680
rect 229 3675 2345 3676
rect 8717 1868 8833 11358
rect 11865 12020 12027 13336
rect 11865 1868 12041 12020
rect 12481 5518 14317 7274
rect 8717 1720 12041 1868
<< via3 >>
rect 5477 15100 8439 19650
rect 8833 1868 11865 13336
<< metal4 >>
rect 71 26932 14451 28248
rect 71 19650 14451 25846
rect 71 15100 5477 19650
rect 8439 15100 14451 19650
rect 71 15044 14451 15100
rect 71 13336 14451 13464
rect 71 9374 8833 13336
rect 11865 9374 14451 13336
rect 14427 8214 14451 9374
rect 71 1868 8833 8214
rect 11865 1868 14451 8214
rect 71 260 14451 1868
<< via4 >>
rect 49 25846 14743 26932
rect 33 8214 8833 9374
rect 8833 8214 11865 9374
rect 11865 8214 14427 9374
<< metal5 >>
rect 25 26932 14767 26956
rect 25 25846 49 26932
rect 14743 25846 14767 26932
rect 25 25822 14767 25846
rect 9 9374 14451 9398
rect 9 8214 33 9374
rect 14427 8214 14451 9374
rect 9 8190 14451 8214
use audiodac_drv_half  audiodac_drv_half_0
timestamp 1644660203
transform 1 0 8677 0 1 35642
box -5906 -21361 6044 -7276
use audiodac_drv_half  audiodac_drv_half_1
timestamp 1644660203
transform 1 0 8677 0 -1 -7276
box -5906 -21361 6044 -7276
use audiodac_drv_latch  audiodac_drv_latch_0
timestamp 1721164599
transform 1 0 1480 0 1 39112
box 1834 -27002 3224 -22840
use audiodac_drv_ls  audiodac_drv_ls_0
timestamp 1724508986
transform 1 0 3778 0 1 31945
box -3728 -20005 -570 -15559
use sky130_fd_pr__pfet_g5v0d10v5_VDASXE  sky130_fd_pr__pfet_g5v0d10v5_VDASXE_0 paramcells
timestamp 1644523392
transform 1 0 1305 0 1 22589
box -1258 -5797 1258 5797
use sky130_fd_pr__pfet_g5v0d10v5_VDASXE  sky130_fd_pr__pfet_g5v0d10v5_VDASXE_1
timestamp 1644523392
transform 1 0 1285 0 1 5797
box -1258 -5797 1258 5797
<< labels >>
rlabel metal3 12481 5518 14317 7274 1 out_p
port 3 n signal output
rlabel metal3 12481 21092 14317 22848 1 out_n
port 4 n signal output
rlabel metal3 8717 1720 12041 12020 1 vss
port 7 n ground input
rlabel metal3 5433 6526 8517 19712 1 vdd
port 5 n power input
rlabel metal1 1 12929 103 15196 1 in_hi
port 6 n signal input
rlabel metal3 70 12329 360 12409 1 in_p
port 1 n signal input
rlabel metal3 70 12509 2750 12589 1 in_n
port 2 n signal input
<< end >>
