magic
tech sky130A
magscale 1 2
timestamp 1644523392
<< nwell >>
rect -1258 -5797 1258 5797
<< mvpmos >>
rect -1000 -5500 1000 5500
<< mvpdiff >>
rect -1058 5488 -1000 5500
rect -1058 -5488 -1046 5488
rect -1012 -5488 -1000 5488
rect -1058 -5500 -1000 -5488
rect 1000 5488 1058 5500
rect 1000 -5488 1012 5488
rect 1046 -5488 1058 5488
rect 1000 -5500 1058 -5488
<< mvpdiffc >>
rect -1046 -5488 -1012 5488
rect 1012 -5488 1046 5488
<< mvnsubdiff >>
rect -1192 5719 1192 5731
rect -1192 5685 -1084 5719
rect 1084 5685 1192 5719
rect -1192 5673 1192 5685
rect -1192 5623 -1134 5673
rect -1192 -5623 -1180 5623
rect -1146 -5623 -1134 5623
rect 1134 5623 1192 5673
rect -1192 -5673 -1134 -5623
rect 1134 -5623 1146 5623
rect 1180 -5623 1192 5623
rect 1134 -5673 1192 -5623
rect -1192 -5685 1192 -5673
rect -1192 -5719 -1084 -5685
rect 1084 -5719 1192 -5685
rect -1192 -5731 1192 -5719
<< mvnsubdiffcont >>
rect -1084 5685 1084 5719
rect -1180 -5623 -1146 5623
rect 1146 -5623 1180 5623
rect -1084 -5719 1084 -5685
<< poly >>
rect -1000 5581 1000 5597
rect -1000 5547 -984 5581
rect 984 5547 1000 5581
rect -1000 5500 1000 5547
rect -1000 -5547 1000 -5500
rect -1000 -5581 -984 -5547
rect 984 -5581 1000 -5547
rect -1000 -5597 1000 -5581
<< polycont >>
rect -984 5547 984 5581
rect -984 -5581 984 -5547
<< locali >>
rect -1180 5685 -1084 5719
rect 1084 5685 1180 5719
rect -1180 5623 -1146 5685
rect 1146 5623 1180 5685
rect -1000 5547 -984 5581
rect 984 5547 1000 5581
rect -1046 5488 -1012 5504
rect -1046 -5504 -1012 -5488
rect 1012 5488 1046 5504
rect 1012 -5504 1046 -5488
rect -1000 -5581 -984 -5547
rect 984 -5581 1000 -5547
rect -1180 -5685 -1146 -5623
rect 1146 -5685 1180 -5623
rect -1180 -5719 -1084 -5685
rect 1084 -5719 1180 -5685
<< viali >>
rect -984 5547 984 5581
rect -1046 -5488 -1012 5488
rect 1012 -5488 1046 5488
rect -984 -5581 984 -5547
<< metal1 >>
rect -996 5581 996 5587
rect -996 5547 -984 5581
rect 984 5547 996 5581
rect -996 5541 996 5547
rect -1052 5488 -1006 5500
rect -1052 -5488 -1046 5488
rect -1012 -5488 -1006 5488
rect -1052 -5500 -1006 -5488
rect 1006 5488 1052 5500
rect 1006 -5488 1012 5488
rect 1046 -5488 1052 5488
rect 1006 -5500 1052 -5488
rect -996 -5547 996 -5541
rect -996 -5581 -984 -5547
rect 984 -5581 996 -5547
rect -996 -5587 996 -5581
<< properties >>
string FIXED_BBOX -1163 -5702 1163 5702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 55 l 10 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
