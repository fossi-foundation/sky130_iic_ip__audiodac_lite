magic
tech sky130A
magscale 1 2
timestamp 1721163516
<< nwell >>
rect -1019 -2415 1019 2415
<< mvpmos >>
rect -761 118 -661 2118
rect -603 118 -503 2118
rect -445 118 -345 2118
rect -287 118 -187 2118
rect -129 118 -29 2118
rect 29 118 129 2118
rect 187 118 287 2118
rect 345 118 445 2118
rect 503 118 603 2118
rect 661 118 761 2118
rect -761 -2118 -661 -118
rect -603 -2118 -503 -118
rect -445 -2118 -345 -118
rect -287 -2118 -187 -118
rect -129 -2118 -29 -118
rect 29 -2118 129 -118
rect 187 -2118 287 -118
rect 345 -2118 445 -118
rect 503 -2118 603 -118
rect 661 -2118 761 -118
<< mvpdiff >>
rect -819 2106 -761 2118
rect -819 130 -807 2106
rect -773 130 -761 2106
rect -819 118 -761 130
rect -661 2106 -603 2118
rect -661 130 -649 2106
rect -615 130 -603 2106
rect -661 118 -603 130
rect -503 2106 -445 2118
rect -503 130 -491 2106
rect -457 130 -445 2106
rect -503 118 -445 130
rect -345 2106 -287 2118
rect -345 130 -333 2106
rect -299 130 -287 2106
rect -345 118 -287 130
rect -187 2106 -129 2118
rect -187 130 -175 2106
rect -141 130 -129 2106
rect -187 118 -129 130
rect -29 2106 29 2118
rect -29 130 -17 2106
rect 17 130 29 2106
rect -29 118 29 130
rect 129 2106 187 2118
rect 129 130 141 2106
rect 175 130 187 2106
rect 129 118 187 130
rect 287 2106 345 2118
rect 287 130 299 2106
rect 333 130 345 2106
rect 287 118 345 130
rect 445 2106 503 2118
rect 445 130 457 2106
rect 491 130 503 2106
rect 445 118 503 130
rect 603 2106 661 2118
rect 603 130 615 2106
rect 649 130 661 2106
rect 603 118 661 130
rect 761 2106 819 2118
rect 761 130 773 2106
rect 807 130 819 2106
rect 761 118 819 130
rect -819 -130 -761 -118
rect -819 -2106 -807 -130
rect -773 -2106 -761 -130
rect -819 -2118 -761 -2106
rect -661 -130 -603 -118
rect -661 -2106 -649 -130
rect -615 -2106 -603 -130
rect -661 -2118 -603 -2106
rect -503 -130 -445 -118
rect -503 -2106 -491 -130
rect -457 -2106 -445 -130
rect -503 -2118 -445 -2106
rect -345 -130 -287 -118
rect -345 -2106 -333 -130
rect -299 -2106 -287 -130
rect -345 -2118 -287 -2106
rect -187 -130 -129 -118
rect -187 -2106 -175 -130
rect -141 -2106 -129 -130
rect -187 -2118 -129 -2106
rect -29 -130 29 -118
rect -29 -2106 -17 -130
rect 17 -2106 29 -130
rect -29 -2118 29 -2106
rect 129 -130 187 -118
rect 129 -2106 141 -130
rect 175 -2106 187 -130
rect 129 -2118 187 -2106
rect 287 -130 345 -118
rect 287 -2106 299 -130
rect 333 -2106 345 -130
rect 287 -2118 345 -2106
rect 445 -130 503 -118
rect 445 -2106 457 -130
rect 491 -2106 503 -130
rect 445 -2118 503 -2106
rect 603 -130 661 -118
rect 603 -2106 615 -130
rect 649 -2106 661 -130
rect 603 -2118 661 -2106
rect 761 -130 819 -118
rect 761 -2106 773 -130
rect 807 -2106 819 -130
rect 761 -2118 819 -2106
<< mvpdiffc >>
rect -807 130 -773 2106
rect -649 130 -615 2106
rect -491 130 -457 2106
rect -333 130 -299 2106
rect -175 130 -141 2106
rect -17 130 17 2106
rect 141 130 175 2106
rect 299 130 333 2106
rect 457 130 491 2106
rect 615 130 649 2106
rect 773 130 807 2106
rect -807 -2106 -773 -130
rect -649 -2106 -615 -130
rect -491 -2106 -457 -130
rect -333 -2106 -299 -130
rect -175 -2106 -141 -130
rect -17 -2106 17 -130
rect 141 -2106 175 -130
rect 299 -2106 333 -130
rect 457 -2106 491 -130
rect 615 -2106 649 -130
rect 773 -2106 807 -130
<< mvnsubdiff >>
rect -953 2337 953 2349
rect -953 2303 -845 2337
rect 845 2303 953 2337
rect -953 2291 953 2303
rect -953 2241 -895 2291
rect -953 -2241 -941 2241
rect -907 -2241 -895 2241
rect 895 2241 953 2291
rect -953 -2291 -895 -2241
rect 895 -2241 907 2241
rect 941 -2241 953 2241
rect 895 -2291 953 -2241
rect -953 -2303 953 -2291
rect -953 -2337 -845 -2303
rect 845 -2337 953 -2303
rect -953 -2349 953 -2337
<< mvnsubdiffcont >>
rect -845 2303 845 2337
rect -941 -2241 -907 2241
rect 907 -2241 941 2241
rect -845 -2337 845 -2303
<< poly >>
rect -761 2199 -661 2215
rect -761 2165 -745 2199
rect -677 2165 -661 2199
rect -761 2118 -661 2165
rect -603 2199 -503 2215
rect -603 2165 -587 2199
rect -519 2165 -503 2199
rect -603 2118 -503 2165
rect -445 2199 -345 2215
rect -445 2165 -429 2199
rect -361 2165 -345 2199
rect -445 2118 -345 2165
rect -287 2199 -187 2215
rect -287 2165 -271 2199
rect -203 2165 -187 2199
rect -287 2118 -187 2165
rect -129 2199 -29 2215
rect -129 2165 -113 2199
rect -45 2165 -29 2199
rect -129 2118 -29 2165
rect 29 2199 129 2215
rect 29 2165 45 2199
rect 113 2165 129 2199
rect 29 2118 129 2165
rect 187 2199 287 2215
rect 187 2165 203 2199
rect 271 2165 287 2199
rect 187 2118 287 2165
rect 345 2199 445 2215
rect 345 2165 361 2199
rect 429 2165 445 2199
rect 345 2118 445 2165
rect 503 2199 603 2215
rect 503 2165 519 2199
rect 587 2165 603 2199
rect 503 2118 603 2165
rect 661 2199 761 2215
rect 661 2165 677 2199
rect 745 2165 761 2199
rect 661 2118 761 2165
rect -761 71 -661 118
rect -761 37 -745 71
rect -677 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -587 71
rect -519 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -429 71
rect -361 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -271 71
rect -203 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -113 71
rect -45 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 45 71
rect 113 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 203 71
rect 271 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 361 71
rect 429 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 519 71
rect 587 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 677 71
rect 745 37 761 71
rect 661 21 761 37
rect -761 -37 -661 -21
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -761 -118 -661 -71
rect -603 -37 -503 -21
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -603 -118 -503 -71
rect -445 -37 -345 -21
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -445 -118 -345 -71
rect -287 -37 -187 -21
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -287 -118 -187 -71
rect -129 -37 -29 -21
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect -129 -118 -29 -71
rect 29 -37 129 -21
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 29 -118 129 -71
rect 187 -37 287 -21
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 187 -118 287 -71
rect 345 -37 445 -21
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 345 -118 445 -71
rect 503 -37 603 -21
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 503 -118 603 -71
rect 661 -37 761 -21
rect 661 -71 677 -37
rect 745 -71 761 -37
rect 661 -118 761 -71
rect -761 -2165 -661 -2118
rect -761 -2199 -745 -2165
rect -677 -2199 -661 -2165
rect -761 -2215 -661 -2199
rect -603 -2165 -503 -2118
rect -603 -2199 -587 -2165
rect -519 -2199 -503 -2165
rect -603 -2215 -503 -2199
rect -445 -2165 -345 -2118
rect -445 -2199 -429 -2165
rect -361 -2199 -345 -2165
rect -445 -2215 -345 -2199
rect -287 -2165 -187 -2118
rect -287 -2199 -271 -2165
rect -203 -2199 -187 -2165
rect -287 -2215 -187 -2199
rect -129 -2165 -29 -2118
rect -129 -2199 -113 -2165
rect -45 -2199 -29 -2165
rect -129 -2215 -29 -2199
rect 29 -2165 129 -2118
rect 29 -2199 45 -2165
rect 113 -2199 129 -2165
rect 29 -2215 129 -2199
rect 187 -2165 287 -2118
rect 187 -2199 203 -2165
rect 271 -2199 287 -2165
rect 187 -2215 287 -2199
rect 345 -2165 445 -2118
rect 345 -2199 361 -2165
rect 429 -2199 445 -2165
rect 345 -2215 445 -2199
rect 503 -2165 603 -2118
rect 503 -2199 519 -2165
rect 587 -2199 603 -2165
rect 503 -2215 603 -2199
rect 661 -2165 761 -2118
rect 661 -2199 677 -2165
rect 745 -2199 761 -2165
rect 661 -2215 761 -2199
<< polycont >>
rect -745 2165 -677 2199
rect -587 2165 -519 2199
rect -429 2165 -361 2199
rect -271 2165 -203 2199
rect -113 2165 -45 2199
rect 45 2165 113 2199
rect 203 2165 271 2199
rect 361 2165 429 2199
rect 519 2165 587 2199
rect 677 2165 745 2199
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect -745 -2199 -677 -2165
rect -587 -2199 -519 -2165
rect -429 -2199 -361 -2165
rect -271 -2199 -203 -2165
rect -113 -2199 -45 -2165
rect 45 -2199 113 -2165
rect 203 -2199 271 -2165
rect 361 -2199 429 -2165
rect 519 -2199 587 -2165
rect 677 -2199 745 -2165
<< locali >>
rect -941 2303 -845 2337
rect 845 2303 941 2337
rect -941 2241 -907 2303
rect 907 2241 941 2303
rect -761 2165 -745 2199
rect -677 2165 -661 2199
rect -603 2165 -587 2199
rect -519 2165 -503 2199
rect -445 2165 -429 2199
rect -361 2165 -345 2199
rect -287 2165 -271 2199
rect -203 2165 -187 2199
rect -129 2165 -113 2199
rect -45 2165 -29 2199
rect 29 2165 45 2199
rect 113 2165 129 2199
rect 187 2165 203 2199
rect 271 2165 287 2199
rect 345 2165 361 2199
rect 429 2165 445 2199
rect 503 2165 519 2199
rect 587 2165 603 2199
rect 661 2165 677 2199
rect 745 2165 761 2199
rect -807 2106 -773 2122
rect -807 114 -773 130
rect -649 2106 -615 2122
rect -649 114 -615 130
rect -491 2106 -457 2122
rect -491 114 -457 130
rect -333 2106 -299 2122
rect -333 114 -299 130
rect -175 2106 -141 2122
rect -175 114 -141 130
rect -17 2106 17 2122
rect -17 114 17 130
rect 141 2106 175 2122
rect 141 114 175 130
rect 299 2106 333 2122
rect 299 114 333 130
rect 457 2106 491 2122
rect 457 114 491 130
rect 615 2106 649 2122
rect 615 114 649 130
rect 773 2106 807 2122
rect 773 114 807 130
rect -761 37 -745 71
rect -677 37 -661 71
rect -603 37 -587 71
rect -519 37 -503 71
rect -445 37 -429 71
rect -361 37 -345 71
rect -287 37 -271 71
rect -203 37 -187 71
rect -129 37 -113 71
rect -45 37 -29 71
rect 29 37 45 71
rect 113 37 129 71
rect 187 37 203 71
rect 271 37 287 71
rect 345 37 361 71
rect 429 37 445 71
rect 503 37 519 71
rect 587 37 603 71
rect 661 37 677 71
rect 745 37 761 71
rect -761 -71 -745 -37
rect -677 -71 -661 -37
rect -603 -71 -587 -37
rect -519 -71 -503 -37
rect -445 -71 -429 -37
rect -361 -71 -345 -37
rect -287 -71 -271 -37
rect -203 -71 -187 -37
rect -129 -71 -113 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 113 -71 129 -37
rect 187 -71 203 -37
rect 271 -71 287 -37
rect 345 -71 361 -37
rect 429 -71 445 -37
rect 503 -71 519 -37
rect 587 -71 603 -37
rect 661 -71 677 -37
rect 745 -71 761 -37
rect -807 -130 -773 -114
rect -807 -2122 -773 -2106
rect -649 -130 -615 -114
rect -649 -2122 -615 -2106
rect -491 -130 -457 -114
rect -491 -2122 -457 -2106
rect -333 -130 -299 -114
rect -333 -2122 -299 -2106
rect -175 -130 -141 -114
rect -175 -2122 -141 -2106
rect -17 -130 17 -114
rect -17 -2122 17 -2106
rect 141 -130 175 -114
rect 141 -2122 175 -2106
rect 299 -130 333 -114
rect 299 -2122 333 -2106
rect 457 -130 491 -114
rect 457 -2122 491 -2106
rect 615 -130 649 -114
rect 615 -2122 649 -2106
rect 773 -130 807 -114
rect 773 -2122 807 -2106
rect -761 -2199 -745 -2165
rect -677 -2199 -661 -2165
rect -603 -2199 -587 -2165
rect -519 -2199 -503 -2165
rect -445 -2199 -429 -2165
rect -361 -2199 -345 -2165
rect -287 -2199 -271 -2165
rect -203 -2199 -187 -2165
rect -129 -2199 -113 -2165
rect -45 -2199 -29 -2165
rect 29 -2199 45 -2165
rect 113 -2199 129 -2165
rect 187 -2199 203 -2165
rect 271 -2199 287 -2165
rect 345 -2199 361 -2165
rect 429 -2199 445 -2165
rect 503 -2199 519 -2165
rect 587 -2199 603 -2165
rect 661 -2199 677 -2165
rect 745 -2199 761 -2165
rect -941 -2303 -907 -2241
rect 907 -2303 941 -2241
rect -941 -2337 -845 -2303
rect 845 -2337 941 -2303
<< viali >>
rect -745 2165 -677 2199
rect -587 2165 -519 2199
rect -429 2165 -361 2199
rect -271 2165 -203 2199
rect -113 2165 -45 2199
rect 45 2165 113 2199
rect 203 2165 271 2199
rect 361 2165 429 2199
rect 519 2165 587 2199
rect 677 2165 745 2199
rect -807 130 -773 2106
rect -649 130 -615 2106
rect -491 130 -457 2106
rect -333 130 -299 2106
rect -175 130 -141 2106
rect -17 130 17 2106
rect 141 130 175 2106
rect 299 130 333 2106
rect 457 130 491 2106
rect 615 130 649 2106
rect 773 130 807 2106
rect -745 37 -677 71
rect -587 37 -519 71
rect -429 37 -361 71
rect -271 37 -203 71
rect -113 37 -45 71
rect 45 37 113 71
rect 203 37 271 71
rect 361 37 429 71
rect 519 37 587 71
rect 677 37 745 71
rect -745 -71 -677 -37
rect -587 -71 -519 -37
rect -429 -71 -361 -37
rect -271 -71 -203 -37
rect -113 -71 -45 -37
rect 45 -71 113 -37
rect 203 -71 271 -37
rect 361 -71 429 -37
rect 519 -71 587 -37
rect 677 -71 745 -37
rect -807 -2106 -773 -130
rect -649 -2106 -615 -130
rect -491 -2106 -457 -130
rect -333 -2106 -299 -130
rect -175 -2106 -141 -130
rect -17 -2106 17 -130
rect 141 -2106 175 -130
rect 299 -2106 333 -130
rect 457 -2106 491 -130
rect 615 -2106 649 -130
rect 773 -2106 807 -130
rect -745 -2199 -677 -2165
rect -587 -2199 -519 -2165
rect -429 -2199 -361 -2165
rect -271 -2199 -203 -2165
rect -113 -2199 -45 -2165
rect 45 -2199 113 -2165
rect 203 -2199 271 -2165
rect 361 -2199 429 -2165
rect 519 -2199 587 -2165
rect 677 -2199 745 -2165
<< metal1 >>
rect -757 2199 -665 2205
rect -757 2165 -745 2199
rect -677 2165 -665 2199
rect -757 2159 -665 2165
rect -599 2199 -507 2205
rect -599 2165 -587 2199
rect -519 2165 -507 2199
rect -599 2159 -507 2165
rect -441 2199 -349 2205
rect -441 2165 -429 2199
rect -361 2165 -349 2199
rect -441 2159 -349 2165
rect -283 2199 -191 2205
rect -283 2165 -271 2199
rect -203 2165 -191 2199
rect -283 2159 -191 2165
rect -125 2199 -33 2205
rect -125 2165 -113 2199
rect -45 2165 -33 2199
rect -125 2159 -33 2165
rect 33 2199 125 2205
rect 33 2165 45 2199
rect 113 2165 125 2199
rect 33 2159 125 2165
rect 191 2199 283 2205
rect 191 2165 203 2199
rect 271 2165 283 2199
rect 191 2159 283 2165
rect 349 2199 441 2205
rect 349 2165 361 2199
rect 429 2165 441 2199
rect 349 2159 441 2165
rect 507 2199 599 2205
rect 507 2165 519 2199
rect 587 2165 599 2199
rect 507 2159 599 2165
rect 665 2199 757 2205
rect 665 2165 677 2199
rect 745 2165 757 2199
rect 665 2159 757 2165
rect -813 2106 -767 2118
rect -813 130 -807 2106
rect -773 130 -767 2106
rect -813 118 -767 130
rect -655 2106 -609 2118
rect -655 130 -649 2106
rect -615 130 -609 2106
rect -655 118 -609 130
rect -497 2106 -451 2118
rect -497 130 -491 2106
rect -457 130 -451 2106
rect -497 118 -451 130
rect -339 2106 -293 2118
rect -339 130 -333 2106
rect -299 130 -293 2106
rect -339 118 -293 130
rect -181 2106 -135 2118
rect -181 130 -175 2106
rect -141 130 -135 2106
rect -181 118 -135 130
rect -23 2106 23 2118
rect -23 130 -17 2106
rect 17 130 23 2106
rect -23 118 23 130
rect 135 2106 181 2118
rect 135 130 141 2106
rect 175 130 181 2106
rect 135 118 181 130
rect 293 2106 339 2118
rect 293 130 299 2106
rect 333 130 339 2106
rect 293 118 339 130
rect 451 2106 497 2118
rect 451 130 457 2106
rect 491 130 497 2106
rect 451 118 497 130
rect 609 2106 655 2118
rect 609 130 615 2106
rect 649 130 655 2106
rect 609 118 655 130
rect 767 2106 813 2118
rect 767 130 773 2106
rect 807 130 813 2106
rect 767 118 813 130
rect -757 71 -665 77
rect -757 37 -745 71
rect -677 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -587 71
rect -519 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -429 71
rect -361 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -271 71
rect -203 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -113 71
rect -45 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 45 71
rect 113 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 203 71
rect 271 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 361 71
rect 429 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 519 71
rect 587 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 677 71
rect 745 37 757 71
rect 665 31 757 37
rect -757 -37 -665 -31
rect -757 -71 -745 -37
rect -677 -71 -665 -37
rect -757 -77 -665 -71
rect -599 -37 -507 -31
rect -599 -71 -587 -37
rect -519 -71 -507 -37
rect -599 -77 -507 -71
rect -441 -37 -349 -31
rect -441 -71 -429 -37
rect -361 -71 -349 -37
rect -441 -77 -349 -71
rect -283 -37 -191 -31
rect -283 -71 -271 -37
rect -203 -71 -191 -37
rect -283 -77 -191 -71
rect -125 -37 -33 -31
rect -125 -71 -113 -37
rect -45 -71 -33 -37
rect -125 -77 -33 -71
rect 33 -37 125 -31
rect 33 -71 45 -37
rect 113 -71 125 -37
rect 33 -77 125 -71
rect 191 -37 283 -31
rect 191 -71 203 -37
rect 271 -71 283 -37
rect 191 -77 283 -71
rect 349 -37 441 -31
rect 349 -71 361 -37
rect 429 -71 441 -37
rect 349 -77 441 -71
rect 507 -37 599 -31
rect 507 -71 519 -37
rect 587 -71 599 -37
rect 507 -77 599 -71
rect 665 -37 757 -31
rect 665 -71 677 -37
rect 745 -71 757 -37
rect 665 -77 757 -71
rect -813 -130 -767 -118
rect -813 -2106 -807 -130
rect -773 -2106 -767 -130
rect -813 -2118 -767 -2106
rect -655 -130 -609 -118
rect -655 -2106 -649 -130
rect -615 -2106 -609 -130
rect -655 -2118 -609 -2106
rect -497 -130 -451 -118
rect -497 -2106 -491 -130
rect -457 -2106 -451 -130
rect -497 -2118 -451 -2106
rect -339 -130 -293 -118
rect -339 -2106 -333 -130
rect -299 -2106 -293 -130
rect -339 -2118 -293 -2106
rect -181 -130 -135 -118
rect -181 -2106 -175 -130
rect -141 -2106 -135 -130
rect -181 -2118 -135 -2106
rect -23 -130 23 -118
rect -23 -2106 -17 -130
rect 17 -2106 23 -130
rect -23 -2118 23 -2106
rect 135 -130 181 -118
rect 135 -2106 141 -130
rect 175 -2106 181 -130
rect 135 -2118 181 -2106
rect 293 -130 339 -118
rect 293 -2106 299 -130
rect 333 -2106 339 -130
rect 293 -2118 339 -2106
rect 451 -130 497 -118
rect 451 -2106 457 -130
rect 491 -2106 497 -130
rect 451 -2118 497 -2106
rect 609 -130 655 -118
rect 609 -2106 615 -130
rect 649 -2106 655 -130
rect 609 -2118 655 -2106
rect 767 -130 813 -118
rect 767 -2106 773 -130
rect 807 -2106 813 -130
rect 767 -2118 813 -2106
rect -757 -2165 -665 -2159
rect -757 -2199 -745 -2165
rect -677 -2199 -665 -2165
rect -757 -2205 -665 -2199
rect -599 -2165 -507 -2159
rect -599 -2199 -587 -2165
rect -519 -2199 -507 -2165
rect -599 -2205 -507 -2199
rect -441 -2165 -349 -2159
rect -441 -2199 -429 -2165
rect -361 -2199 -349 -2165
rect -441 -2205 -349 -2199
rect -283 -2165 -191 -2159
rect -283 -2199 -271 -2165
rect -203 -2199 -191 -2165
rect -283 -2205 -191 -2199
rect -125 -2165 -33 -2159
rect -125 -2199 -113 -2165
rect -45 -2199 -33 -2165
rect -125 -2205 -33 -2199
rect 33 -2165 125 -2159
rect 33 -2199 45 -2165
rect 113 -2199 125 -2165
rect 33 -2205 125 -2199
rect 191 -2165 283 -2159
rect 191 -2199 203 -2165
rect 271 -2199 283 -2165
rect 191 -2205 283 -2199
rect 349 -2165 441 -2159
rect 349 -2199 361 -2165
rect 429 -2199 441 -2165
rect 349 -2205 441 -2199
rect 507 -2165 599 -2159
rect 507 -2199 519 -2165
rect 587 -2199 599 -2165
rect 507 -2205 599 -2199
rect 665 -2165 757 -2159
rect 665 -2199 677 -2165
rect 745 -2199 757 -2165
rect 665 -2205 757 -2199
<< properties >>
string FIXED_BBOX -924 -2320 924 2320
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 0.5 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
