magic
tech sky130A
magscale 1 2
timestamp 1721164599
<< nwell >>
rect 1834 -25434 3224 -22840
<< pwell >>
rect 1864 -27002 3194 -25486
<< mvnmos >>
rect 2092 -26744 2192 -25744
rect 2250 -26744 2350 -25744
rect 2708 -26744 2808 -25744
rect 2866 -26744 2966 -25744
<< mvpmos >>
rect 2092 -25138 2192 -23138
rect 2250 -25138 2350 -23138
rect 2708 -25138 2808 -23138
rect 2866 -25138 2966 -23138
<< mvndiff >>
rect 2034 -25756 2092 -25744
rect 2034 -26732 2046 -25756
rect 2080 -26732 2092 -25756
rect 2034 -26744 2092 -26732
rect 2192 -25756 2250 -25744
rect 2192 -26732 2204 -25756
rect 2238 -26732 2250 -25756
rect 2192 -26744 2250 -26732
rect 2350 -25756 2408 -25744
rect 2350 -26732 2362 -25756
rect 2396 -26732 2408 -25756
rect 2350 -26744 2408 -26732
rect 2650 -25756 2708 -25744
rect 2650 -26732 2662 -25756
rect 2696 -26732 2708 -25756
rect 2650 -26744 2708 -26732
rect 2808 -25756 2866 -25744
rect 2808 -26732 2820 -25756
rect 2854 -26732 2866 -25756
rect 2808 -26744 2866 -26732
rect 2966 -25756 3024 -25744
rect 2966 -26732 2978 -25756
rect 3012 -26732 3024 -25756
rect 2966 -26744 3024 -26732
<< mvpdiff >>
rect 2034 -23150 2092 -23138
rect 2034 -25126 2046 -23150
rect 2080 -25126 2092 -23150
rect 2034 -25138 2092 -25126
rect 2192 -23150 2250 -23138
rect 2192 -25126 2204 -23150
rect 2238 -25126 2250 -23150
rect 2192 -25138 2250 -25126
rect 2350 -23150 2408 -23138
rect 2350 -25126 2362 -23150
rect 2396 -25126 2408 -23150
rect 2350 -25138 2408 -25126
rect 2650 -23150 2708 -23138
rect 2650 -25126 2662 -23150
rect 2696 -25126 2708 -23150
rect 2650 -25138 2708 -25126
rect 2808 -23150 2866 -23138
rect 2808 -25126 2820 -23150
rect 2854 -25126 2866 -23150
rect 2808 -25138 2866 -25126
rect 2966 -23150 3024 -23138
rect 2966 -25126 2978 -23150
rect 3012 -25126 3024 -23150
rect 2966 -25138 3024 -25126
<< mvndiffc >>
rect 2046 -26732 2080 -25756
rect 2204 -26732 2238 -25756
rect 2362 -26732 2396 -25756
rect 2662 -26732 2696 -25756
rect 2820 -26732 2854 -25756
rect 2978 -26732 3012 -25756
<< mvpdiffc >>
rect 2046 -25126 2080 -23150
rect 2204 -25126 2238 -23150
rect 2362 -25126 2396 -23150
rect 2662 -25126 2696 -23150
rect 2820 -25126 2854 -23150
rect 2978 -25126 3012 -23150
<< mvpsubdiff >>
rect 1900 -25534 3158 -25522
rect 1900 -25568 2008 -25534
rect 2434 -25568 2624 -25534
rect 3050 -25568 3158 -25534
rect 1900 -25580 3158 -25568
rect 1900 -25630 1958 -25580
rect 1900 -26858 1912 -25630
rect 1946 -26858 1958 -25630
rect 2484 -25630 2574 -25580
rect 1900 -26908 1958 -26858
rect 2484 -26858 2496 -25630
rect 2562 -26858 2574 -25630
rect 3100 -25630 3158 -25580
rect 2484 -26908 2574 -26858
rect 3100 -26858 3112 -25630
rect 3146 -26858 3158 -25630
rect 3100 -26908 3158 -26858
rect 1900 -26920 3158 -26908
rect 1900 -26954 2008 -26920
rect 2434 -26954 2624 -26920
rect 3050 -26954 3158 -26920
rect 1900 -26966 3158 -26954
<< mvnsubdiff >>
rect 1900 -22918 3158 -22906
rect 1900 -22952 2008 -22918
rect 2434 -22952 2624 -22918
rect 3050 -22952 3158 -22918
rect 1900 -22964 3158 -22952
rect 1900 -23014 1958 -22964
rect 1900 -25260 1912 -23014
rect 1946 -25260 1958 -23014
rect 2484 -23014 2574 -22964
rect 1900 -25310 1958 -25260
rect 2484 -25260 2496 -23014
rect 2562 -25260 2574 -23014
rect 3100 -23014 3158 -22964
rect 2484 -25310 2574 -25260
rect 3100 -25260 3112 -23014
rect 3146 -25260 3158 -23014
rect 3100 -25310 3158 -25260
rect 1900 -25322 3158 -25310
rect 1900 -25356 2008 -25322
rect 2434 -25356 2624 -25322
rect 3050 -25356 3158 -25322
rect 1900 -25368 3158 -25356
<< mvpsubdiffcont >>
rect 2008 -25568 2434 -25534
rect 2624 -25568 3050 -25534
rect 1912 -26858 1946 -25630
rect 2496 -26858 2562 -25630
rect 3112 -26858 3146 -25630
rect 2008 -26954 2434 -26920
rect 2624 -26954 3050 -26920
<< mvnsubdiffcont >>
rect 2008 -22952 2434 -22918
rect 2624 -22952 3050 -22918
rect 1912 -25260 1946 -23014
rect 2496 -25260 2562 -23014
rect 3112 -25260 3146 -23014
rect 2008 -25356 2434 -25322
rect 2624 -25356 3050 -25322
<< poly >>
rect 2092 -23056 2192 -23040
rect 2092 -23090 2108 -23056
rect 2176 -23090 2192 -23056
rect 2092 -23138 2192 -23090
rect 2250 -23056 2350 -23040
rect 2250 -23090 2266 -23056
rect 2334 -23090 2350 -23056
rect 2250 -23138 2350 -23090
rect 2092 -25186 2192 -25138
rect 2092 -25220 2108 -25186
rect 2176 -25220 2192 -25186
rect 2092 -25236 2192 -25220
rect 2250 -25186 2350 -25138
rect 2250 -25220 2266 -25186
rect 2334 -25220 2350 -25186
rect 2250 -25236 2350 -25220
rect 2708 -23056 2808 -23040
rect 2708 -23090 2724 -23056
rect 2792 -23090 2808 -23056
rect 2708 -23138 2808 -23090
rect 2866 -23056 2966 -23040
rect 2866 -23090 2882 -23056
rect 2950 -23090 2966 -23056
rect 2866 -23138 2966 -23090
rect 2708 -25186 2808 -25138
rect 2708 -25220 2724 -25186
rect 2792 -25220 2808 -25186
rect 2708 -25236 2808 -25220
rect 2866 -25186 2966 -25138
rect 2866 -25220 2882 -25186
rect 2950 -25220 2966 -25186
rect 2866 -25236 2966 -25220
rect 2092 -25672 2192 -25656
rect 2092 -25706 2108 -25672
rect 2176 -25706 2192 -25672
rect 2092 -25744 2192 -25706
rect 2250 -25672 2350 -25656
rect 2250 -25706 2266 -25672
rect 2334 -25706 2350 -25672
rect 2250 -25744 2350 -25706
rect 2092 -26782 2192 -26744
rect 2092 -26816 2108 -26782
rect 2176 -26816 2192 -26782
rect 2092 -26832 2192 -26816
rect 2250 -26782 2350 -26744
rect 2250 -26816 2266 -26782
rect 2334 -26816 2350 -26782
rect 2250 -26832 2350 -26816
rect 2708 -25672 2808 -25656
rect 2708 -25706 2724 -25672
rect 2792 -25706 2808 -25672
rect 2708 -25744 2808 -25706
rect 2866 -25672 2966 -25656
rect 2866 -25706 2882 -25672
rect 2950 -25706 2966 -25672
rect 2866 -25744 2966 -25706
rect 2708 -26782 2808 -26744
rect 2708 -26816 2724 -26782
rect 2792 -26816 2808 -26782
rect 2708 -26832 2808 -26816
rect 2866 -26782 2966 -26744
rect 2866 -26816 2882 -26782
rect 2950 -26816 2966 -26782
rect 2866 -26832 2966 -26816
<< polycont >>
rect 2108 -23090 2176 -23056
rect 2266 -23090 2334 -23056
rect 2108 -25220 2176 -25186
rect 2266 -25220 2334 -25186
rect 2724 -23090 2792 -23056
rect 2882 -23090 2950 -23056
rect 2724 -25220 2792 -25186
rect 2882 -25220 2950 -25186
rect 2108 -25706 2176 -25672
rect 2266 -25706 2334 -25672
rect 2108 -26816 2176 -26782
rect 2266 -26816 2334 -26782
rect 2724 -25706 2792 -25672
rect 2882 -25706 2950 -25672
rect 2724 -26816 2792 -26782
rect 2882 -26816 2950 -26782
<< locali >>
rect 1912 -22952 2008 -22918
rect 2434 -22952 2624 -22918
rect 3050 -22952 3146 -22918
rect 1912 -23014 1946 -22952
rect 2496 -23014 2562 -22952
rect 2092 -23090 2108 -23056
rect 2176 -23090 2192 -23056
rect 2250 -23090 2266 -23056
rect 2334 -23090 2350 -23056
rect 2046 -23150 2080 -23134
rect 2046 -25142 2080 -25126
rect 2204 -23150 2238 -23134
rect 2204 -25142 2238 -25126
rect 2362 -23150 2396 -23134
rect 3112 -23014 3146 -22952
rect 2708 -23090 2724 -23056
rect 2792 -23090 2808 -23056
rect 2866 -23090 2882 -23056
rect 2950 -23090 2966 -23056
rect 2662 -23150 2696 -23134
rect 2362 -25142 2396 -25126
rect 2092 -25220 2108 -25186
rect 2176 -25220 2192 -25186
rect 2250 -25220 2266 -25186
rect 2334 -25220 2350 -25186
rect 1912 -25322 1946 -25260
rect 2662 -25142 2696 -25126
rect 2820 -23150 2854 -23134
rect 2820 -25142 2854 -25126
rect 2978 -23150 3012 -23134
rect 2978 -25142 3012 -25126
rect 2708 -25220 2724 -25186
rect 2792 -25220 2808 -25186
rect 2866 -25220 2882 -25186
rect 2950 -25220 2966 -25186
rect 2496 -25322 2562 -25260
rect 3112 -25322 3146 -25260
rect 1912 -25356 2008 -25322
rect 2434 -25356 2624 -25322
rect 3050 -25356 3146 -25322
rect 1912 -25568 2008 -25534
rect 2434 -25568 2624 -25534
rect 3050 -25568 3146 -25534
rect 1912 -25630 1946 -25568
rect 2496 -25630 2562 -25568
rect 2092 -25706 2108 -25672
rect 2176 -25706 2192 -25672
rect 2250 -25706 2266 -25672
rect 2334 -25706 2350 -25672
rect 2046 -25756 2080 -25740
rect 2046 -26748 2080 -26732
rect 2204 -25756 2238 -25740
rect 2204 -26748 2238 -26732
rect 2362 -25756 2396 -25740
rect 3112 -25630 3146 -25568
rect 2708 -25706 2724 -25672
rect 2792 -25706 2808 -25672
rect 2866 -25706 2882 -25672
rect 2950 -25706 2966 -25672
rect 2662 -25756 2696 -25740
rect 2362 -26748 2396 -26732
rect 2092 -26816 2108 -26782
rect 2176 -26816 2192 -26782
rect 2250 -26816 2266 -26782
rect 2334 -26816 2350 -26782
rect 1912 -26920 1946 -26858
rect 2662 -26748 2696 -26732
rect 2820 -25756 2854 -25740
rect 2820 -26748 2854 -26732
rect 2978 -25756 3012 -25740
rect 2978 -26748 3012 -26732
rect 2708 -26816 2724 -26782
rect 2792 -26816 2808 -26782
rect 2866 -26816 2882 -26782
rect 2950 -26816 2966 -26782
rect 2496 -26920 2562 -26858
rect 3112 -26920 3146 -26858
rect 1912 -26954 2008 -26920
rect 2434 -26954 2624 -26920
rect 3050 -26954 3146 -26920
<< viali >>
rect 2108 -23090 2176 -23056
rect 2266 -23090 2334 -23056
rect 2046 -25126 2080 -23150
rect 2204 -25126 2238 -23150
rect 2362 -25126 2396 -23150
rect 2724 -23090 2792 -23056
rect 2882 -23090 2950 -23056
rect 2488 -23322 2496 -23152
rect 2496 -23322 2562 -23152
rect 2562 -23322 2572 -23152
rect 2108 -25220 2176 -25186
rect 2266 -25220 2334 -25186
rect 2662 -25126 2696 -23150
rect 2820 -25126 2854 -23150
rect 2978 -25126 3012 -23150
rect 2724 -25220 2792 -25186
rect 2882 -25220 2950 -25186
rect 2108 -25706 2176 -25672
rect 2266 -25706 2334 -25672
rect 2046 -26732 2080 -25756
rect 2204 -26732 2238 -25756
rect 2362 -26732 2396 -25756
rect 2724 -25706 2792 -25672
rect 2882 -25706 2950 -25672
rect 2486 -26706 2496 -26536
rect 2496 -26706 2562 -26536
rect 2562 -26706 2570 -26536
rect 2108 -26816 2176 -26782
rect 2266 -26816 2334 -26782
rect 2662 -26732 2696 -25756
rect 2820 -26732 2854 -25756
rect 2978 -26732 3012 -25756
rect 2724 -26816 2792 -26782
rect 2882 -26816 2950 -26782
<< metal1 >>
rect 2090 -23055 2346 -23046
rect 1947 -23056 2349 -23055
rect 1947 -23090 2108 -23056
rect 2176 -23090 2266 -23056
rect 2334 -23090 2349 -23056
rect 2703 -23056 3117 -23041
rect 2703 -23087 2724 -23056
rect 1947 -23101 2349 -23090
rect 2710 -23090 2724 -23087
rect 2792 -23090 2882 -23056
rect 2950 -23087 3117 -23056
rect 2950 -23090 2966 -23087
rect 2710 -23092 2966 -23090
rect 2712 -23096 2804 -23092
rect 2870 -23096 2962 -23092
rect 1947 -25180 1993 -23101
rect 2040 -23150 2086 -23138
rect 2040 -23152 2046 -23150
rect 2080 -23152 2086 -23150
rect 2198 -23150 2244 -23138
rect 2028 -23322 2038 -23152
rect 2090 -23322 2100 -23152
rect 2040 -25126 2046 -23322
rect 2080 -25126 2086 -23322
rect 2198 -25018 2204 -23150
rect 2238 -25018 2244 -23150
rect 2356 -23150 2402 -23138
rect 2356 -23152 2362 -23150
rect 2396 -23152 2402 -23150
rect 2482 -23152 2578 -23140
rect 2656 -23150 2702 -23138
rect 2656 -23152 2662 -23150
rect 2696 -23152 2702 -23150
rect 2814 -23150 2860 -23138
rect 2344 -23322 2354 -23152
rect 2406 -23322 2416 -23152
rect 2478 -23322 2488 -23152
rect 2572 -23322 2582 -23152
rect 2644 -23322 2654 -23152
rect 2706 -23322 2716 -23152
rect 2180 -25116 2190 -25018
rect 2256 -25116 2266 -25018
rect 2040 -25138 2086 -25126
rect 2198 -25126 2204 -25116
rect 2238 -25126 2244 -25116
rect 2198 -25138 2244 -25126
rect 2356 -25126 2362 -23322
rect 2396 -25126 2402 -23322
rect 2482 -23334 2578 -23322
rect 2356 -25138 2402 -25126
rect 2656 -25126 2662 -23322
rect 2696 -25126 2702 -23322
rect 2814 -25018 2820 -23150
rect 2854 -25018 2860 -23150
rect 2972 -23150 3018 -23138
rect 2972 -23152 2978 -23150
rect 3012 -23152 3018 -23150
rect 2960 -23322 2970 -23152
rect 3022 -23322 3032 -23152
rect 2794 -25116 2804 -25018
rect 2870 -25116 2880 -25018
rect 2656 -25138 2702 -25126
rect 2814 -25126 2820 -25116
rect 2854 -25126 2860 -25116
rect 2814 -25138 2860 -25126
rect 2972 -25126 2978 -23322
rect 3012 -25126 3018 -23322
rect 2972 -25138 3018 -25126
rect 1947 -25186 2348 -25180
rect 2712 -25184 2964 -25180
rect 3071 -25184 3117 -23087
rect 1947 -25220 2108 -25186
rect 2176 -25220 2266 -25186
rect 2334 -25220 2348 -25186
rect 1947 -25226 2348 -25220
rect 2096 -25516 2348 -25226
rect 2702 -25186 3117 -25184
rect 2702 -25220 2724 -25186
rect 2792 -25220 2882 -25186
rect 2950 -25220 3117 -25186
rect 2702 -25230 3117 -25220
rect 2480 -25302 2578 -25296
rect 2712 -25302 2964 -25230
rect 2578 -25368 2964 -25302
rect 2480 -25374 2578 -25368
rect 2480 -25516 2578 -25510
rect 2096 -25582 2480 -25516
rect 2096 -25664 2348 -25582
rect 2480 -25588 2578 -25582
rect 2712 -25650 2964 -25368
rect 1924 -25672 2348 -25664
rect 1924 -25706 2108 -25672
rect 2176 -25706 2266 -25672
rect 2334 -25706 2348 -25672
rect 2700 -25672 3114 -25650
rect 2700 -25702 2724 -25672
rect 1924 -25712 2348 -25706
rect 2712 -25706 2724 -25702
rect 2792 -25706 2882 -25672
rect 2950 -25702 3114 -25672
rect 2950 -25706 2964 -25702
rect 2712 -25712 2964 -25706
rect 1924 -26782 1976 -25712
rect 2040 -25756 2086 -25744
rect 2040 -26536 2046 -25756
rect 2080 -26536 2086 -25756
rect 2180 -25838 2190 -25740
rect 2256 -25838 2266 -25740
rect 2356 -25756 2402 -25744
rect 2028 -26706 2038 -26536
rect 2090 -26706 2100 -26536
rect 2040 -26732 2046 -26706
rect 2080 -26732 2086 -26706
rect 2040 -26744 2086 -26732
rect 2198 -26732 2204 -25838
rect 2238 -26732 2244 -25838
rect 2356 -26536 2362 -25756
rect 2396 -26536 2402 -25756
rect 2656 -25756 2702 -25744
rect 2480 -26536 2576 -26524
rect 2656 -26536 2662 -25756
rect 2696 -26536 2702 -25756
rect 2794 -25838 2804 -25740
rect 2870 -25838 2880 -25740
rect 2972 -25756 3018 -25744
rect 2344 -26706 2354 -26536
rect 2406 -26706 2416 -26536
rect 2476 -26706 2486 -26536
rect 2570 -26706 2580 -26536
rect 2644 -26706 2654 -26536
rect 2706 -26706 2716 -26536
rect 2198 -26744 2244 -26732
rect 2356 -26732 2362 -26706
rect 2396 -26732 2402 -26706
rect 2480 -26718 2576 -26706
rect 2356 -26744 2402 -26732
rect 2656 -26732 2662 -26706
rect 2696 -26732 2702 -26706
rect 2656 -26744 2702 -26732
rect 2814 -26732 2820 -25838
rect 2854 -26732 2860 -25838
rect 2972 -26536 2978 -25756
rect 3012 -26536 3018 -25756
rect 2958 -26706 2968 -26536
rect 3020 -26706 3030 -26536
rect 2814 -26744 2860 -26732
rect 2972 -26732 2978 -26706
rect 3012 -26732 3018 -26706
rect 2972 -26744 3018 -26732
rect 2096 -26780 2188 -26776
rect 2254 -26780 2346 -26776
rect 2712 -26778 2804 -26776
rect 2870 -26778 2962 -26776
rect 2094 -26782 2350 -26780
rect 1924 -26816 2108 -26782
rect 2176 -26816 2266 -26782
rect 2334 -26816 2350 -26782
rect 1924 -26824 2350 -26816
rect 2708 -26782 2964 -26778
rect 2708 -26816 2724 -26782
rect 2792 -26816 2882 -26782
rect 2950 -26786 2964 -26782
rect 3062 -26786 3114 -25702
rect 2950 -26816 3114 -26786
rect 1924 -26834 2344 -26824
rect 2708 -26838 3114 -26816
<< via1 >>
rect 2038 -23322 2046 -23152
rect 2046 -23322 2080 -23152
rect 2080 -23322 2090 -23152
rect 2354 -23322 2362 -23152
rect 2362 -23322 2396 -23152
rect 2396 -23322 2406 -23152
rect 2488 -23322 2572 -23152
rect 2654 -23322 2662 -23152
rect 2662 -23322 2696 -23152
rect 2696 -23322 2706 -23152
rect 2190 -25116 2204 -25018
rect 2204 -25116 2238 -25018
rect 2238 -25116 2256 -25018
rect 2970 -23322 2978 -23152
rect 2978 -23322 3012 -23152
rect 3012 -23322 3022 -23152
rect 2804 -25116 2820 -25018
rect 2820 -25116 2854 -25018
rect 2854 -25116 2870 -25018
rect 2480 -25368 2578 -25302
rect 2480 -25582 2578 -25516
rect 2190 -25756 2256 -25740
rect 2190 -25838 2204 -25756
rect 2204 -25838 2238 -25756
rect 2238 -25838 2256 -25756
rect 2038 -26706 2046 -26536
rect 2046 -26706 2080 -26536
rect 2080 -26706 2090 -26536
rect 2804 -25756 2870 -25740
rect 2804 -25838 2820 -25756
rect 2820 -25838 2854 -25756
rect 2854 -25838 2870 -25756
rect 2354 -26706 2362 -26536
rect 2362 -26706 2396 -26536
rect 2396 -26706 2406 -26536
rect 2486 -26706 2570 -26536
rect 2654 -26706 2662 -26536
rect 2662 -26706 2696 -26536
rect 2696 -26706 2706 -26536
rect 2968 -26706 2978 -26536
rect 2978 -26706 3012 -26536
rect 3012 -26706 3020 -26536
<< metal2 >>
rect 2038 -23152 2090 -23142
rect 2354 -23152 2406 -23142
rect 2488 -23152 2572 -23142
rect 2654 -23152 2706 -23142
rect 2970 -23152 3022 -23142
rect 2090 -23322 2354 -23152
rect 2406 -23322 2488 -23152
rect 2572 -23322 2654 -23152
rect 2706 -23322 2970 -23152
rect 2038 -23332 2090 -23322
rect 2354 -23332 2406 -23322
rect 2488 -23332 2572 -23322
rect 2654 -23332 2706 -23322
rect 2970 -23332 3022 -23322
rect 2190 -25018 2256 -25008
rect 2190 -25302 2256 -25116
rect 2804 -25018 2870 -25008
rect 2190 -25368 2480 -25302
rect 2578 -25368 2584 -25302
rect 2190 -25740 2256 -25368
rect 2804 -25516 2870 -25116
rect 2474 -25582 2480 -25516
rect 2578 -25582 2870 -25516
rect 2190 -25848 2256 -25838
rect 2804 -25740 2870 -25582
rect 2804 -25848 2870 -25838
rect 2038 -26536 2090 -26526
rect 2354 -26536 2406 -26526
rect 2486 -26536 2570 -26526
rect 2654 -26536 2706 -26526
rect 2968 -26536 3020 -26526
rect 2090 -26706 2354 -26536
rect 2406 -26706 2486 -26536
rect 2570 -26706 2654 -26536
rect 2706 -26706 2968 -26536
rect 2038 -26716 2090 -26706
rect 2354 -26716 2406 -26706
rect 2486 -26716 2570 -26706
rect 2654 -26716 2706 -26706
rect 2968 -26716 3020 -26706
<< labels >>
rlabel metal2 2804 -25740 2870 -25116 1 in_n
port 2 n
rlabel metal2 2190 -25740 2256 -25116 1 in_p
port 1 n
rlabel metal2 2090 -26706 2354 -26536 1 vss
port 4 n
rlabel metal2 2090 -23322 2354 -23152 1 vdd_hi
port 3 n
<< end >>
