magic
tech sky130A
timestamp 1644523392
<< nwell >>
rect -312 -248 312 248
<< mvpmos >>
rect -183 -100 -133 100
rect -104 -100 -54 100
rect -25 -100 25 100
rect 54 -100 104 100
rect 133 -100 183 100
<< mvpdiff >>
rect -212 94 -183 100
rect -212 -94 -206 94
rect -189 -94 -183 94
rect -212 -100 -183 -94
rect -133 94 -104 100
rect -133 -94 -127 94
rect -110 -94 -104 94
rect -133 -100 -104 -94
rect -54 94 -25 100
rect -54 -94 -48 94
rect -31 -94 -25 94
rect -54 -100 -25 -94
rect 25 94 54 100
rect 25 -94 31 94
rect 48 -94 54 94
rect 25 -100 54 -94
rect 104 94 133 100
rect 104 -94 110 94
rect 127 -94 133 94
rect 104 -100 133 -94
rect 183 94 212 100
rect 183 -94 189 94
rect 206 -94 212 94
rect 183 -100 212 -94
<< mvpdiffc >>
rect -206 -94 -189 94
rect -127 -94 -110 94
rect -48 -94 -31 94
rect 31 -94 48 94
rect 110 -94 127 94
rect 189 -94 206 94
<< mvnsubdiff >>
rect -279 209 279 215
rect -279 192 -225 209
rect 225 192 279 209
rect -279 186 279 192
rect -279 161 -250 186
rect -279 -161 -273 161
rect -256 -161 -250 161
rect 250 161 279 186
rect -279 -186 -250 -161
rect 250 -161 256 161
rect 273 -161 279 161
rect 250 -186 279 -161
rect -279 -192 279 -186
rect -279 -209 -225 -192
rect 225 -209 279 -192
rect -279 -215 279 -209
<< mvnsubdiffcont >>
rect -225 192 225 209
rect -273 -161 -256 161
rect 256 -161 273 161
rect -225 -209 225 -192
<< poly >>
rect -183 141 -133 149
rect -183 124 -175 141
rect -141 124 -133 141
rect -183 100 -133 124
rect -104 141 -54 149
rect -104 124 -96 141
rect -62 124 -54 141
rect -104 100 -54 124
rect -25 141 25 149
rect -25 124 -17 141
rect 17 124 25 141
rect -25 100 25 124
rect 54 141 104 149
rect 54 124 62 141
rect 96 124 104 141
rect 54 100 104 124
rect 133 141 183 149
rect 133 124 141 141
rect 175 124 183 141
rect 133 100 183 124
rect -183 -124 -133 -100
rect -183 -141 -175 -124
rect -141 -141 -133 -124
rect -183 -149 -133 -141
rect -104 -124 -54 -100
rect -104 -141 -96 -124
rect -62 -141 -54 -124
rect -104 -149 -54 -141
rect -25 -124 25 -100
rect -25 -141 -17 -124
rect 17 -141 25 -124
rect -25 -149 25 -141
rect 54 -124 104 -100
rect 54 -141 62 -124
rect 96 -141 104 -124
rect 54 -149 104 -141
rect 133 -124 183 -100
rect 133 -141 141 -124
rect 175 -141 183 -124
rect 133 -149 183 -141
<< polycont >>
rect -175 124 -141 141
rect -96 124 -62 141
rect -17 124 17 141
rect 62 124 96 141
rect 141 124 175 141
rect -175 -141 -141 -124
rect -96 -141 -62 -124
rect -17 -141 17 -124
rect 62 -141 96 -124
rect 141 -141 175 -124
<< locali >>
rect -273 192 -225 209
rect 225 192 273 209
rect -273 161 -256 192
rect 256 161 273 192
rect -183 124 -175 141
rect -141 124 -133 141
rect -104 124 -96 141
rect -62 124 -54 141
rect -25 124 -17 141
rect 17 124 25 141
rect 54 124 62 141
rect 96 124 104 141
rect 133 124 141 141
rect 175 124 183 141
rect -206 94 -189 102
rect -206 -102 -189 -94
rect -127 94 -110 102
rect -127 -102 -110 -94
rect -48 94 -31 102
rect -48 -102 -31 -94
rect 31 94 48 102
rect 31 -102 48 -94
rect 110 94 127 102
rect 110 -102 127 -94
rect 189 94 206 102
rect 189 -102 206 -94
rect -183 -141 -175 -124
rect -141 -141 -133 -124
rect -104 -141 -96 -124
rect -62 -141 -54 -124
rect -25 -141 -17 -124
rect 17 -141 25 -124
rect 54 -141 62 -124
rect 96 -141 104 -124
rect 133 -141 141 -124
rect 175 -141 183 -124
rect -273 -192 -256 -161
rect 256 -192 273 -161
rect -273 -209 -225 -192
rect 225 -209 273 -192
<< viali >>
rect -175 124 -141 141
rect -96 124 -62 141
rect -17 124 17 141
rect 62 124 96 141
rect 141 124 175 141
rect -206 -94 -189 94
rect -127 -94 -110 94
rect -48 -94 -31 94
rect 31 -94 48 94
rect 110 -94 127 94
rect 189 -94 206 94
rect -175 -141 -141 -124
rect -96 -141 -62 -124
rect -17 -141 17 -124
rect 62 -141 96 -124
rect 141 -141 175 -124
<< metal1 >>
rect -181 141 -135 144
rect -181 124 -175 141
rect -141 124 -135 141
rect -181 121 -135 124
rect -102 141 -56 144
rect -102 124 -96 141
rect -62 124 -56 141
rect -102 121 -56 124
rect -23 141 23 144
rect -23 124 -17 141
rect 17 124 23 141
rect -23 121 23 124
rect 56 141 102 144
rect 56 124 62 141
rect 96 124 102 141
rect 56 121 102 124
rect 135 141 181 144
rect 135 124 141 141
rect 175 124 181 141
rect 135 121 181 124
rect -209 94 -186 100
rect -209 -94 -206 94
rect -189 -94 -186 94
rect -209 -100 -186 -94
rect -130 94 -107 100
rect -130 -94 -127 94
rect -110 -94 -107 94
rect -130 -100 -107 -94
rect -51 94 -28 100
rect -51 -94 -48 94
rect -31 -94 -28 94
rect -51 -100 -28 -94
rect 28 94 51 100
rect 28 -94 31 94
rect 48 -94 51 94
rect 28 -100 51 -94
rect 107 94 130 100
rect 107 -94 110 94
rect 127 -94 130 94
rect 107 -100 130 -94
rect 186 94 209 100
rect 186 -94 189 94
rect 206 -94 209 94
rect 186 -100 209 -94
rect -181 -124 -135 -121
rect -181 -141 -175 -124
rect -141 -141 -135 -124
rect -181 -144 -135 -141
rect -102 -124 -56 -121
rect -102 -141 -96 -124
rect -62 -141 -56 -124
rect -102 -144 -56 -141
rect -23 -124 23 -121
rect -23 -141 -17 -124
rect 17 -141 23 -124
rect -23 -144 23 -141
rect 56 -124 102 -121
rect 56 -141 62 -124
rect 96 -141 102 -124
rect 56 -144 102 -141
rect 135 -124 181 -121
rect 135 -141 141 -124
rect 175 -141 181 -124
rect 135 -144 181 -141
<< properties >>
string FIXED_BBOX -264 -201 264 201
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
