magic
tech sky130A
timestamp 1644523392
<< pwell >>
rect -397 -629 397 629
<< mvnnmos >>
rect -283 -500 -193 500
rect -164 -500 -74 500
rect -45 -500 45 500
rect 74 -500 164 500
rect 193 -500 283 500
<< mvndiff >>
rect -312 494 -283 500
rect -312 -494 -306 494
rect -289 -494 -283 494
rect -312 -500 -283 -494
rect -193 494 -164 500
rect -193 -494 -187 494
rect -170 -494 -164 494
rect -193 -500 -164 -494
rect -74 494 -45 500
rect -74 -494 -68 494
rect -51 -494 -45 494
rect -74 -500 -45 -494
rect 45 494 74 500
rect 45 -494 51 494
rect 68 -494 74 494
rect 45 -500 74 -494
rect 164 494 193 500
rect 164 -494 170 494
rect 187 -494 193 494
rect 164 -500 193 -494
rect 283 494 312 500
rect 283 -494 289 494
rect 306 -494 312 494
rect 283 -500 312 -494
<< mvndiffc >>
rect -306 -494 -289 494
rect -187 -494 -170 494
rect -68 -494 -51 494
rect 51 -494 68 494
rect 170 -494 187 494
rect 289 -494 306 494
<< mvpsubdiff >>
rect -379 605 379 611
rect -379 588 -325 605
rect 325 588 379 605
rect -379 582 379 588
rect -379 557 -350 582
rect -379 -557 -373 557
rect -356 -557 -350 557
rect 350 557 379 582
rect -379 -582 -350 -557
rect 350 -557 356 557
rect 373 -557 379 557
rect 350 -582 379 -557
rect -379 -588 379 -582
rect -379 -605 -325 -588
rect 325 -605 379 -588
rect -379 -611 379 -605
<< mvpsubdiffcont >>
rect -325 588 325 605
rect -373 -557 -356 557
rect 356 -557 373 557
rect -325 -605 325 -588
<< poly >>
rect -283 536 -193 544
rect -283 519 -275 536
rect -201 519 -193 536
rect -283 500 -193 519
rect -164 536 -74 544
rect -164 519 -156 536
rect -82 519 -74 536
rect -164 500 -74 519
rect -45 536 45 544
rect -45 519 -37 536
rect 37 519 45 536
rect -45 500 45 519
rect 74 536 164 544
rect 74 519 82 536
rect 156 519 164 536
rect 74 500 164 519
rect 193 536 283 544
rect 193 519 201 536
rect 275 519 283 536
rect 193 500 283 519
rect -283 -519 -193 -500
rect -283 -536 -275 -519
rect -201 -536 -193 -519
rect -283 -544 -193 -536
rect -164 -519 -74 -500
rect -164 -536 -156 -519
rect -82 -536 -74 -519
rect -164 -544 -74 -536
rect -45 -519 45 -500
rect -45 -536 -37 -519
rect 37 -536 45 -519
rect -45 -544 45 -536
rect 74 -519 164 -500
rect 74 -536 82 -519
rect 156 -536 164 -519
rect 74 -544 164 -536
rect 193 -519 283 -500
rect 193 -536 201 -519
rect 275 -536 283 -519
rect 193 -544 283 -536
<< polycont >>
rect -275 519 -201 536
rect -156 519 -82 536
rect -37 519 37 536
rect 82 519 156 536
rect 201 519 275 536
rect -275 -536 -201 -519
rect -156 -536 -82 -519
rect -37 -536 37 -519
rect 82 -536 156 -519
rect 201 -536 275 -519
<< locali >>
rect -373 588 -325 605
rect 325 588 373 605
rect -373 557 -356 588
rect 356 557 373 588
rect -283 519 -275 536
rect -201 519 -193 536
rect -164 519 -156 536
rect -82 519 -74 536
rect -45 519 -37 536
rect 37 519 45 536
rect 74 519 82 536
rect 156 519 164 536
rect 193 519 201 536
rect 275 519 283 536
rect -306 494 -289 502
rect -306 -502 -289 -494
rect -187 494 -170 502
rect -187 -502 -170 -494
rect -68 494 -51 502
rect -68 -502 -51 -494
rect 51 494 68 502
rect 51 -502 68 -494
rect 170 494 187 502
rect 170 -502 187 -494
rect 289 494 306 502
rect 289 -502 306 -494
rect -283 -536 -275 -519
rect -201 -536 -193 -519
rect -164 -536 -156 -519
rect -82 -536 -74 -519
rect -45 -536 -37 -519
rect 37 -536 45 -519
rect 74 -536 82 -519
rect 156 -536 164 -519
rect 193 -536 201 -519
rect 275 -536 283 -519
rect -373 -588 -356 -557
rect 356 -588 373 -557
rect -373 -605 -325 -588
rect 325 -605 373 -588
<< viali >>
rect -275 519 -201 536
rect -156 519 -82 536
rect -37 519 37 536
rect 82 519 156 536
rect 201 519 275 536
rect -306 -494 -289 494
rect -187 -494 -170 494
rect -68 -494 -51 494
rect 51 -494 68 494
rect 170 -494 187 494
rect 289 -494 306 494
rect -275 -536 -201 -519
rect -156 -536 -82 -519
rect -37 -536 37 -519
rect 82 -536 156 -519
rect 201 -536 275 -519
<< metal1 >>
rect -281 536 -195 539
rect -281 519 -275 536
rect -201 519 -195 536
rect -281 516 -195 519
rect -162 536 -76 539
rect -162 519 -156 536
rect -82 519 -76 536
rect -162 516 -76 519
rect -43 536 43 539
rect -43 519 -37 536
rect 37 519 43 536
rect -43 516 43 519
rect 76 536 162 539
rect 76 519 82 536
rect 156 519 162 536
rect 76 516 162 519
rect 195 536 281 539
rect 195 519 201 536
rect 275 519 281 536
rect 195 516 281 519
rect -309 494 -286 500
rect -309 -494 -306 494
rect -289 -494 -286 494
rect -309 -500 -286 -494
rect -190 494 -167 500
rect -190 -494 -187 494
rect -170 -494 -167 494
rect -190 -500 -167 -494
rect -71 494 -48 500
rect -71 -494 -68 494
rect -51 -494 -48 494
rect -71 -500 -48 -494
rect 48 494 71 500
rect 48 -494 51 494
rect 68 -494 71 494
rect 48 -500 71 -494
rect 167 494 190 500
rect 167 -494 170 494
rect 187 -494 190 494
rect 167 -500 190 -494
rect 286 494 309 500
rect 286 -494 289 494
rect 306 -494 309 494
rect 286 -500 309 -494
rect -281 -519 -195 -516
rect -281 -536 -275 -519
rect -201 -536 -195 -519
rect -281 -539 -195 -536
rect -162 -519 -76 -516
rect -162 -536 -156 -519
rect -82 -536 -76 -519
rect -162 -539 -76 -536
rect -43 -519 43 -516
rect -43 -536 -37 -519
rect 37 -536 43 -519
rect -43 -539 43 -536
rect 76 -519 162 -516
rect 76 -536 82 -519
rect 156 -536 162 -519
rect 76 -539 162 -536
rect 195 -519 281 -516
rect 195 -536 201 -519
rect 275 -536 281 -519
rect 195 -539 281 -536
<< properties >>
string FIXED_BBOX -364 -596 364 596
string gencell sky130_fd_pr__nfet_05v0_nvt
string library sky130
string parameters w 10 l 0.90 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.90 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
