magic
tech sky130A
magscale 1 2
timestamp 1721163516
<< pwell >>
rect -989 -1258 989 1258
<< mvnmos >>
rect -761 -1000 -661 1000
rect -603 -1000 -503 1000
rect -445 -1000 -345 1000
rect -287 -1000 -187 1000
rect -129 -1000 -29 1000
rect 29 -1000 129 1000
rect 187 -1000 287 1000
rect 345 -1000 445 1000
rect 503 -1000 603 1000
rect 661 -1000 761 1000
<< mvndiff >>
rect -819 988 -761 1000
rect -819 -988 -807 988
rect -773 -988 -761 988
rect -819 -1000 -761 -988
rect -661 988 -603 1000
rect -661 -988 -649 988
rect -615 -988 -603 988
rect -661 -1000 -603 -988
rect -503 988 -445 1000
rect -503 -988 -491 988
rect -457 -988 -445 988
rect -503 -1000 -445 -988
rect -345 988 -287 1000
rect -345 -988 -333 988
rect -299 -988 -287 988
rect -345 -1000 -287 -988
rect -187 988 -129 1000
rect -187 -988 -175 988
rect -141 -988 -129 988
rect -187 -1000 -129 -988
rect -29 988 29 1000
rect -29 -988 -17 988
rect 17 -988 29 988
rect -29 -1000 29 -988
rect 129 988 187 1000
rect 129 -988 141 988
rect 175 -988 187 988
rect 129 -1000 187 -988
rect 287 988 345 1000
rect 287 -988 299 988
rect 333 -988 345 988
rect 287 -1000 345 -988
rect 445 988 503 1000
rect 445 -988 457 988
rect 491 -988 503 988
rect 445 -1000 503 -988
rect 603 988 661 1000
rect 603 -988 615 988
rect 649 -988 661 988
rect 603 -1000 661 -988
rect 761 988 819 1000
rect 761 -988 773 988
rect 807 -988 819 988
rect 761 -1000 819 -988
<< mvndiffc >>
rect -807 -988 -773 988
rect -649 -988 -615 988
rect -491 -988 -457 988
rect -333 -988 -299 988
rect -175 -988 -141 988
rect -17 -988 17 988
rect 141 -988 175 988
rect 299 -988 333 988
rect 457 -988 491 988
rect 615 -988 649 988
rect 773 -988 807 988
<< mvpsubdiff >>
rect -953 1210 953 1222
rect -953 1176 -845 1210
rect 845 1176 953 1210
rect -953 1164 953 1176
rect -953 1114 -895 1164
rect -953 -1114 -941 1114
rect -907 -1114 -895 1114
rect 895 1114 953 1164
rect -953 -1164 -895 -1114
rect 895 -1114 907 1114
rect 941 -1114 953 1114
rect 895 -1164 953 -1114
rect -953 -1176 953 -1164
rect -953 -1210 -845 -1176
rect 845 -1210 953 -1176
rect -953 -1222 953 -1210
<< mvpsubdiffcont >>
rect -845 1176 845 1210
rect -941 -1114 -907 1114
rect 907 -1114 941 1114
rect -845 -1210 845 -1176
<< poly >>
rect -761 1072 -661 1088
rect -761 1038 -745 1072
rect -677 1038 -661 1072
rect -761 1000 -661 1038
rect -603 1072 -503 1088
rect -603 1038 -587 1072
rect -519 1038 -503 1072
rect -603 1000 -503 1038
rect -445 1072 -345 1088
rect -445 1038 -429 1072
rect -361 1038 -345 1072
rect -445 1000 -345 1038
rect -287 1072 -187 1088
rect -287 1038 -271 1072
rect -203 1038 -187 1072
rect -287 1000 -187 1038
rect -129 1072 -29 1088
rect -129 1038 -113 1072
rect -45 1038 -29 1072
rect -129 1000 -29 1038
rect 29 1072 129 1088
rect 29 1038 45 1072
rect 113 1038 129 1072
rect 29 1000 129 1038
rect 187 1072 287 1088
rect 187 1038 203 1072
rect 271 1038 287 1072
rect 187 1000 287 1038
rect 345 1072 445 1088
rect 345 1038 361 1072
rect 429 1038 445 1072
rect 345 1000 445 1038
rect 503 1072 603 1088
rect 503 1038 519 1072
rect 587 1038 603 1072
rect 503 1000 603 1038
rect 661 1072 761 1088
rect 661 1038 677 1072
rect 745 1038 761 1072
rect 661 1000 761 1038
rect -761 -1038 -661 -1000
rect -761 -1072 -745 -1038
rect -677 -1072 -661 -1038
rect -761 -1088 -661 -1072
rect -603 -1038 -503 -1000
rect -603 -1072 -587 -1038
rect -519 -1072 -503 -1038
rect -603 -1088 -503 -1072
rect -445 -1038 -345 -1000
rect -445 -1072 -429 -1038
rect -361 -1072 -345 -1038
rect -445 -1088 -345 -1072
rect -287 -1038 -187 -1000
rect -287 -1072 -271 -1038
rect -203 -1072 -187 -1038
rect -287 -1088 -187 -1072
rect -129 -1038 -29 -1000
rect -129 -1072 -113 -1038
rect -45 -1072 -29 -1038
rect -129 -1088 -29 -1072
rect 29 -1038 129 -1000
rect 29 -1072 45 -1038
rect 113 -1072 129 -1038
rect 29 -1088 129 -1072
rect 187 -1038 287 -1000
rect 187 -1072 203 -1038
rect 271 -1072 287 -1038
rect 187 -1088 287 -1072
rect 345 -1038 445 -1000
rect 345 -1072 361 -1038
rect 429 -1072 445 -1038
rect 345 -1088 445 -1072
rect 503 -1038 603 -1000
rect 503 -1072 519 -1038
rect 587 -1072 603 -1038
rect 503 -1088 603 -1072
rect 661 -1038 761 -1000
rect 661 -1072 677 -1038
rect 745 -1072 761 -1038
rect 661 -1088 761 -1072
<< polycont >>
rect -745 1038 -677 1072
rect -587 1038 -519 1072
rect -429 1038 -361 1072
rect -271 1038 -203 1072
rect -113 1038 -45 1072
rect 45 1038 113 1072
rect 203 1038 271 1072
rect 361 1038 429 1072
rect 519 1038 587 1072
rect 677 1038 745 1072
rect -745 -1072 -677 -1038
rect -587 -1072 -519 -1038
rect -429 -1072 -361 -1038
rect -271 -1072 -203 -1038
rect -113 -1072 -45 -1038
rect 45 -1072 113 -1038
rect 203 -1072 271 -1038
rect 361 -1072 429 -1038
rect 519 -1072 587 -1038
rect 677 -1072 745 -1038
<< locali >>
rect -941 1176 -845 1210
rect 845 1176 941 1210
rect -941 1114 -907 1176
rect 907 1114 941 1176
rect -761 1038 -745 1072
rect -677 1038 -661 1072
rect -603 1038 -587 1072
rect -519 1038 -503 1072
rect -445 1038 -429 1072
rect -361 1038 -345 1072
rect -287 1038 -271 1072
rect -203 1038 -187 1072
rect -129 1038 -113 1072
rect -45 1038 -29 1072
rect 29 1038 45 1072
rect 113 1038 129 1072
rect 187 1038 203 1072
rect 271 1038 287 1072
rect 345 1038 361 1072
rect 429 1038 445 1072
rect 503 1038 519 1072
rect 587 1038 603 1072
rect 661 1038 677 1072
rect 745 1038 761 1072
rect -807 988 -773 1004
rect -807 -1004 -773 -988
rect -649 988 -615 1004
rect -649 -1004 -615 -988
rect -491 988 -457 1004
rect -491 -1004 -457 -988
rect -333 988 -299 1004
rect -333 -1004 -299 -988
rect -175 988 -141 1004
rect -175 -1004 -141 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 141 988 175 1004
rect 141 -1004 175 -988
rect 299 988 333 1004
rect 299 -1004 333 -988
rect 457 988 491 1004
rect 457 -1004 491 -988
rect 615 988 649 1004
rect 615 -1004 649 -988
rect 773 988 807 1004
rect 773 -1004 807 -988
rect -761 -1072 -745 -1038
rect -677 -1072 -661 -1038
rect -603 -1072 -587 -1038
rect -519 -1072 -503 -1038
rect -445 -1072 -429 -1038
rect -361 -1072 -345 -1038
rect -287 -1072 -271 -1038
rect -203 -1072 -187 -1038
rect -129 -1072 -113 -1038
rect -45 -1072 -29 -1038
rect 29 -1072 45 -1038
rect 113 -1072 129 -1038
rect 187 -1072 203 -1038
rect 271 -1072 287 -1038
rect 345 -1072 361 -1038
rect 429 -1072 445 -1038
rect 503 -1072 519 -1038
rect 587 -1072 603 -1038
rect 661 -1072 677 -1038
rect 745 -1072 761 -1038
rect -941 -1176 -907 -1114
rect 907 -1176 941 -1114
rect -941 -1210 -845 -1176
rect 845 -1210 941 -1176
<< viali >>
rect -745 1038 -677 1072
rect -587 1038 -519 1072
rect -429 1038 -361 1072
rect -271 1038 -203 1072
rect -113 1038 -45 1072
rect 45 1038 113 1072
rect 203 1038 271 1072
rect 361 1038 429 1072
rect 519 1038 587 1072
rect 677 1038 745 1072
rect -807 -988 -773 988
rect -649 -988 -615 988
rect -491 -988 -457 988
rect -333 -988 -299 988
rect -175 -988 -141 988
rect -17 -988 17 988
rect 141 -988 175 988
rect 299 -988 333 988
rect 457 -988 491 988
rect 615 -988 649 988
rect 773 -988 807 988
rect -745 -1072 -677 -1038
rect -587 -1072 -519 -1038
rect -429 -1072 -361 -1038
rect -271 -1072 -203 -1038
rect -113 -1072 -45 -1038
rect 45 -1072 113 -1038
rect 203 -1072 271 -1038
rect 361 -1072 429 -1038
rect 519 -1072 587 -1038
rect 677 -1072 745 -1038
<< metal1 >>
rect -757 1072 -665 1078
rect -757 1038 -745 1072
rect -677 1038 -665 1072
rect -757 1032 -665 1038
rect -599 1072 -507 1078
rect -599 1038 -587 1072
rect -519 1038 -507 1072
rect -599 1032 -507 1038
rect -441 1072 -349 1078
rect -441 1038 -429 1072
rect -361 1038 -349 1072
rect -441 1032 -349 1038
rect -283 1072 -191 1078
rect -283 1038 -271 1072
rect -203 1038 -191 1072
rect -283 1032 -191 1038
rect -125 1072 -33 1078
rect -125 1038 -113 1072
rect -45 1038 -33 1072
rect -125 1032 -33 1038
rect 33 1072 125 1078
rect 33 1038 45 1072
rect 113 1038 125 1072
rect 33 1032 125 1038
rect 191 1072 283 1078
rect 191 1038 203 1072
rect 271 1038 283 1072
rect 191 1032 283 1038
rect 349 1072 441 1078
rect 349 1038 361 1072
rect 429 1038 441 1072
rect 349 1032 441 1038
rect 507 1072 599 1078
rect 507 1038 519 1072
rect 587 1038 599 1072
rect 507 1032 599 1038
rect 665 1072 757 1078
rect 665 1038 677 1072
rect 745 1038 757 1072
rect 665 1032 757 1038
rect -813 988 -767 1000
rect -813 -988 -807 988
rect -773 -988 -767 988
rect -813 -1000 -767 -988
rect -655 988 -609 1000
rect -655 -988 -649 988
rect -615 -988 -609 988
rect -655 -1000 -609 -988
rect -497 988 -451 1000
rect -497 -988 -491 988
rect -457 -988 -451 988
rect -497 -1000 -451 -988
rect -339 988 -293 1000
rect -339 -988 -333 988
rect -299 -988 -293 988
rect -339 -1000 -293 -988
rect -181 988 -135 1000
rect -181 -988 -175 988
rect -141 -988 -135 988
rect -181 -1000 -135 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 135 988 181 1000
rect 135 -988 141 988
rect 175 -988 181 988
rect 135 -1000 181 -988
rect 293 988 339 1000
rect 293 -988 299 988
rect 333 -988 339 988
rect 293 -1000 339 -988
rect 451 988 497 1000
rect 451 -988 457 988
rect 491 -988 497 988
rect 451 -1000 497 -988
rect 609 988 655 1000
rect 609 -988 615 988
rect 649 -988 655 988
rect 609 -1000 655 -988
rect 767 988 813 1000
rect 767 -988 773 988
rect 807 -988 813 988
rect 767 -1000 813 -988
rect -757 -1038 -665 -1032
rect -757 -1072 -745 -1038
rect -677 -1072 -665 -1038
rect -757 -1078 -665 -1072
rect -599 -1038 -507 -1032
rect -599 -1072 -587 -1038
rect -519 -1072 -507 -1038
rect -599 -1078 -507 -1072
rect -441 -1038 -349 -1032
rect -441 -1072 -429 -1038
rect -361 -1072 -349 -1038
rect -441 -1078 -349 -1072
rect -283 -1038 -191 -1032
rect -283 -1072 -271 -1038
rect -203 -1072 -191 -1038
rect -283 -1078 -191 -1072
rect -125 -1038 -33 -1032
rect -125 -1072 -113 -1038
rect -45 -1072 -33 -1038
rect -125 -1078 -33 -1072
rect 33 -1038 125 -1032
rect 33 -1072 45 -1038
rect 113 -1072 125 -1038
rect 33 -1078 125 -1072
rect 191 -1038 283 -1032
rect 191 -1072 203 -1038
rect 271 -1072 283 -1038
rect 191 -1078 283 -1072
rect 349 -1038 441 -1032
rect 349 -1072 361 -1038
rect 429 -1072 441 -1038
rect 349 -1078 441 -1072
rect 507 -1038 599 -1032
rect 507 -1072 519 -1038
rect 587 -1072 599 -1038
rect 507 -1078 599 -1072
rect 665 -1038 757 -1032
rect 665 -1072 677 -1038
rect 745 -1072 757 -1038
rect 665 -1078 757 -1072
<< properties >>
string FIXED_BBOX -924 -1193 924 1193
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 10.0 l 0.5 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
