magic
tech sky130A
timestamp 1644523392
<< nwell >>
rect -509 -1207 509 1207
<< mvpmos >>
rect -380 59 -330 1059
rect -301 59 -251 1059
rect -222 59 -172 1059
rect -143 59 -93 1059
rect -64 59 -14 1059
rect 15 59 65 1059
rect 94 59 144 1059
rect 173 59 223 1059
rect 252 59 302 1059
rect 331 59 381 1059
rect -380 -1059 -330 -59
rect -301 -1059 -251 -59
rect -222 -1059 -172 -59
rect -143 -1059 -93 -59
rect -64 -1059 -14 -59
rect 15 -1059 65 -59
rect 94 -1059 144 -59
rect 173 -1059 223 -59
rect 252 -1059 302 -59
rect 331 -1059 381 -59
<< mvpdiff >>
rect -409 1053 -380 1059
rect -409 65 -403 1053
rect -386 65 -380 1053
rect -409 59 -380 65
rect -330 1053 -301 1059
rect -330 65 -324 1053
rect -307 65 -301 1053
rect -330 59 -301 65
rect -251 1053 -222 1059
rect -251 65 -245 1053
rect -228 65 -222 1053
rect -251 59 -222 65
rect -172 1053 -143 1059
rect -172 65 -166 1053
rect -149 65 -143 1053
rect -172 59 -143 65
rect -93 1053 -64 1059
rect -93 65 -87 1053
rect -70 65 -64 1053
rect -93 59 -64 65
rect -14 1053 15 1059
rect -14 65 -8 1053
rect 9 65 15 1053
rect -14 59 15 65
rect 65 1053 94 1059
rect 65 65 71 1053
rect 88 65 94 1053
rect 65 59 94 65
rect 144 1053 173 1059
rect 144 65 150 1053
rect 167 65 173 1053
rect 144 59 173 65
rect 223 1053 252 1059
rect 223 65 229 1053
rect 246 65 252 1053
rect 223 59 252 65
rect 302 1053 331 1059
rect 302 65 308 1053
rect 325 65 331 1053
rect 302 59 331 65
rect 381 1053 410 1059
rect 381 65 387 1053
rect 404 65 410 1053
rect 381 59 410 65
rect -409 -65 -380 -59
rect -409 -1053 -403 -65
rect -386 -1053 -380 -65
rect -409 -1059 -380 -1053
rect -330 -65 -301 -59
rect -330 -1053 -324 -65
rect -307 -1053 -301 -65
rect -330 -1059 -301 -1053
rect -251 -65 -222 -59
rect -251 -1053 -245 -65
rect -228 -1053 -222 -65
rect -251 -1059 -222 -1053
rect -172 -65 -143 -59
rect -172 -1053 -166 -65
rect -149 -1053 -143 -65
rect -172 -1059 -143 -1053
rect -93 -65 -64 -59
rect -93 -1053 -87 -65
rect -70 -1053 -64 -65
rect -93 -1059 -64 -1053
rect -14 -65 15 -59
rect -14 -1053 -8 -65
rect 9 -1053 15 -65
rect -14 -1059 15 -1053
rect 65 -65 94 -59
rect 65 -1053 71 -65
rect 88 -1053 94 -65
rect 65 -1059 94 -1053
rect 144 -65 173 -59
rect 144 -1053 150 -65
rect 167 -1053 173 -65
rect 144 -1059 173 -1053
rect 223 -65 252 -59
rect 223 -1053 229 -65
rect 246 -1053 252 -65
rect 223 -1059 252 -1053
rect 302 -65 331 -59
rect 302 -1053 308 -65
rect 325 -1053 331 -65
rect 302 -1059 331 -1053
rect 381 -65 410 -59
rect 381 -1053 387 -65
rect 404 -1053 410 -65
rect 381 -1059 410 -1053
<< mvpdiffc >>
rect -403 65 -386 1053
rect -324 65 -307 1053
rect -245 65 -228 1053
rect -166 65 -149 1053
rect -87 65 -70 1053
rect -8 65 9 1053
rect 71 65 88 1053
rect 150 65 167 1053
rect 229 65 246 1053
rect 308 65 325 1053
rect 387 65 404 1053
rect -403 -1053 -386 -65
rect -324 -1053 -307 -65
rect -245 -1053 -228 -65
rect -166 -1053 -149 -65
rect -87 -1053 -70 -65
rect -8 -1053 9 -65
rect 71 -1053 88 -65
rect 150 -1053 167 -65
rect 229 -1053 246 -65
rect 308 -1053 325 -65
rect 387 -1053 404 -65
<< mvnsubdiff >>
rect -476 1168 476 1174
rect -476 1151 -422 1168
rect 422 1151 476 1168
rect -476 1145 476 1151
rect -476 1120 -447 1145
rect -476 -1120 -470 1120
rect -453 -1120 -447 1120
rect 447 1120 476 1145
rect -476 -1145 -447 -1120
rect 447 -1120 453 1120
rect 470 -1120 476 1120
rect 447 -1145 476 -1120
rect -476 -1151 476 -1145
rect -476 -1168 -422 -1151
rect 422 -1168 476 -1151
rect -476 -1174 476 -1168
<< mvnsubdiffcont >>
rect -422 1151 422 1168
rect -470 -1120 -453 1120
rect 453 -1120 470 1120
rect -422 -1168 422 -1151
<< poly >>
rect -380 1100 -330 1108
rect -380 1083 -372 1100
rect -338 1083 -330 1100
rect -380 1059 -330 1083
rect -301 1100 -251 1108
rect -301 1083 -293 1100
rect -259 1083 -251 1100
rect -301 1059 -251 1083
rect -222 1100 -172 1108
rect -222 1083 -214 1100
rect -180 1083 -172 1100
rect -222 1059 -172 1083
rect -143 1100 -93 1108
rect -143 1083 -135 1100
rect -101 1083 -93 1100
rect -143 1059 -93 1083
rect -64 1100 -14 1108
rect -64 1083 -56 1100
rect -22 1083 -14 1100
rect -64 1059 -14 1083
rect 15 1100 65 1108
rect 15 1083 23 1100
rect 57 1083 65 1100
rect 15 1059 65 1083
rect 94 1100 144 1108
rect 94 1083 102 1100
rect 136 1083 144 1100
rect 94 1059 144 1083
rect 173 1100 223 1108
rect 173 1083 181 1100
rect 215 1083 223 1100
rect 173 1059 223 1083
rect 252 1100 302 1108
rect 252 1083 260 1100
rect 294 1083 302 1100
rect 252 1059 302 1083
rect 331 1100 381 1108
rect 331 1083 339 1100
rect 373 1083 381 1100
rect 331 1059 381 1083
rect -380 35 -330 59
rect -380 18 -372 35
rect -338 18 -330 35
rect -380 -18 -330 18
rect -380 -35 -372 -18
rect -338 -35 -330 -18
rect -380 -59 -330 -35
rect -301 35 -251 59
rect -301 18 -293 35
rect -259 18 -251 35
rect -301 -18 -251 18
rect -301 -35 -293 -18
rect -259 -35 -251 -18
rect -301 -59 -251 -35
rect -222 35 -172 59
rect -222 18 -214 35
rect -180 18 -172 35
rect -222 -18 -172 18
rect -222 -35 -214 -18
rect -180 -35 -172 -18
rect -222 -59 -172 -35
rect -143 35 -93 59
rect -143 18 -135 35
rect -101 18 -93 35
rect -143 -18 -93 18
rect -143 -35 -135 -18
rect -101 -35 -93 -18
rect -143 -59 -93 -35
rect -64 35 -14 59
rect -64 18 -56 35
rect -22 18 -14 35
rect -64 -18 -14 18
rect -64 -35 -56 -18
rect -22 -35 -14 -18
rect -64 -59 -14 -35
rect 15 35 65 59
rect 15 18 23 35
rect 57 18 65 35
rect 15 -18 65 18
rect 15 -35 23 -18
rect 57 -35 65 -18
rect 15 -59 65 -35
rect 94 35 144 59
rect 94 18 102 35
rect 136 18 144 35
rect 94 -18 144 18
rect 94 -35 102 -18
rect 136 -35 144 -18
rect 94 -59 144 -35
rect 173 35 223 59
rect 173 18 181 35
rect 215 18 223 35
rect 173 -18 223 18
rect 173 -35 181 -18
rect 215 -35 223 -18
rect 173 -59 223 -35
rect 252 35 302 59
rect 252 18 260 35
rect 294 18 302 35
rect 252 -18 302 18
rect 252 -35 260 -18
rect 294 -35 302 -18
rect 252 -59 302 -35
rect 331 35 381 59
rect 331 18 339 35
rect 373 18 381 35
rect 331 -18 381 18
rect 331 -35 339 -18
rect 373 -35 381 -18
rect 331 -59 381 -35
rect -380 -1083 -330 -1059
rect -380 -1100 -372 -1083
rect -338 -1100 -330 -1083
rect -380 -1108 -330 -1100
rect -301 -1083 -251 -1059
rect -301 -1100 -293 -1083
rect -259 -1100 -251 -1083
rect -301 -1108 -251 -1100
rect -222 -1083 -172 -1059
rect -222 -1100 -214 -1083
rect -180 -1100 -172 -1083
rect -222 -1108 -172 -1100
rect -143 -1083 -93 -1059
rect -143 -1100 -135 -1083
rect -101 -1100 -93 -1083
rect -143 -1108 -93 -1100
rect -64 -1083 -14 -1059
rect -64 -1100 -56 -1083
rect -22 -1100 -14 -1083
rect -64 -1108 -14 -1100
rect 15 -1083 65 -1059
rect 15 -1100 23 -1083
rect 57 -1100 65 -1083
rect 15 -1108 65 -1100
rect 94 -1083 144 -1059
rect 94 -1100 102 -1083
rect 136 -1100 144 -1083
rect 94 -1108 144 -1100
rect 173 -1083 223 -1059
rect 173 -1100 181 -1083
rect 215 -1100 223 -1083
rect 173 -1108 223 -1100
rect 252 -1083 302 -1059
rect 252 -1100 260 -1083
rect 294 -1100 302 -1083
rect 252 -1108 302 -1100
rect 331 -1083 381 -1059
rect 331 -1100 339 -1083
rect 373 -1100 381 -1083
rect 331 -1108 381 -1100
<< polycont >>
rect -372 1083 -338 1100
rect -293 1083 -259 1100
rect -214 1083 -180 1100
rect -135 1083 -101 1100
rect -56 1083 -22 1100
rect 23 1083 57 1100
rect 102 1083 136 1100
rect 181 1083 215 1100
rect 260 1083 294 1100
rect 339 1083 373 1100
rect -372 18 -338 35
rect -372 -35 -338 -18
rect -293 18 -259 35
rect -293 -35 -259 -18
rect -214 18 -180 35
rect -214 -35 -180 -18
rect -135 18 -101 35
rect -135 -35 -101 -18
rect -56 18 -22 35
rect -56 -35 -22 -18
rect 23 18 57 35
rect 23 -35 57 -18
rect 102 18 136 35
rect 102 -35 136 -18
rect 181 18 215 35
rect 181 -35 215 -18
rect 260 18 294 35
rect 260 -35 294 -18
rect 339 18 373 35
rect 339 -35 373 -18
rect -372 -1100 -338 -1083
rect -293 -1100 -259 -1083
rect -214 -1100 -180 -1083
rect -135 -1100 -101 -1083
rect -56 -1100 -22 -1083
rect 23 -1100 57 -1083
rect 102 -1100 136 -1083
rect 181 -1100 215 -1083
rect 260 -1100 294 -1083
rect 339 -1100 373 -1083
<< locali >>
rect -470 1151 -422 1168
rect 422 1151 470 1168
rect -470 1120 -453 1151
rect 453 1120 470 1151
rect -380 1083 -372 1100
rect -338 1083 -330 1100
rect -301 1083 -293 1100
rect -259 1083 -251 1100
rect -222 1083 -214 1100
rect -180 1083 -172 1100
rect -143 1083 -135 1100
rect -101 1083 -93 1100
rect -64 1083 -56 1100
rect -22 1083 -14 1100
rect 15 1083 23 1100
rect 57 1083 65 1100
rect 94 1083 102 1100
rect 136 1083 144 1100
rect 173 1083 181 1100
rect 215 1083 223 1100
rect 252 1083 260 1100
rect 294 1083 302 1100
rect 331 1083 339 1100
rect 373 1083 381 1100
rect -403 1053 -386 1061
rect -403 57 -386 65
rect -324 1053 -307 1061
rect -324 57 -307 65
rect -245 1053 -228 1061
rect -245 57 -228 65
rect -166 1053 -149 1061
rect -166 57 -149 65
rect -87 1053 -70 1061
rect -87 57 -70 65
rect -8 1053 9 1061
rect -8 57 9 65
rect 71 1053 88 1061
rect 71 57 88 65
rect 150 1053 167 1061
rect 150 57 167 65
rect 229 1053 246 1061
rect 229 57 246 65
rect 308 1053 325 1061
rect 308 57 325 65
rect 387 1053 404 1061
rect 387 57 404 65
rect -380 18 -372 35
rect -338 18 -330 35
rect -301 18 -293 35
rect -259 18 -251 35
rect -222 18 -214 35
rect -180 18 -172 35
rect -143 18 -135 35
rect -101 18 -93 35
rect -64 18 -56 35
rect -22 18 -14 35
rect 15 18 23 35
rect 57 18 65 35
rect 94 18 102 35
rect 136 18 144 35
rect 173 18 181 35
rect 215 18 223 35
rect 252 18 260 35
rect 294 18 302 35
rect 331 18 339 35
rect 373 18 381 35
rect -380 -35 -372 -18
rect -338 -35 -330 -18
rect -301 -35 -293 -18
rect -259 -35 -251 -18
rect -222 -35 -214 -18
rect -180 -35 -172 -18
rect -143 -35 -135 -18
rect -101 -35 -93 -18
rect -64 -35 -56 -18
rect -22 -35 -14 -18
rect 15 -35 23 -18
rect 57 -35 65 -18
rect 94 -35 102 -18
rect 136 -35 144 -18
rect 173 -35 181 -18
rect 215 -35 223 -18
rect 252 -35 260 -18
rect 294 -35 302 -18
rect 331 -35 339 -18
rect 373 -35 381 -18
rect -403 -65 -386 -57
rect -403 -1061 -386 -1053
rect -324 -65 -307 -57
rect -324 -1061 -307 -1053
rect -245 -65 -228 -57
rect -245 -1061 -228 -1053
rect -166 -65 -149 -57
rect -166 -1061 -149 -1053
rect -87 -65 -70 -57
rect -87 -1061 -70 -1053
rect -8 -65 9 -57
rect -8 -1061 9 -1053
rect 71 -65 88 -57
rect 71 -1061 88 -1053
rect 150 -65 167 -57
rect 150 -1061 167 -1053
rect 229 -65 246 -57
rect 229 -1061 246 -1053
rect 308 -65 325 -57
rect 308 -1061 325 -1053
rect 387 -65 404 -57
rect 387 -1061 404 -1053
rect -380 -1100 -372 -1083
rect -338 -1100 -330 -1083
rect -301 -1100 -293 -1083
rect -259 -1100 -251 -1083
rect -222 -1100 -214 -1083
rect -180 -1100 -172 -1083
rect -143 -1100 -135 -1083
rect -101 -1100 -93 -1083
rect -64 -1100 -56 -1083
rect -22 -1100 -14 -1083
rect 15 -1100 23 -1083
rect 57 -1100 65 -1083
rect 94 -1100 102 -1083
rect 136 -1100 144 -1083
rect 173 -1100 181 -1083
rect 215 -1100 223 -1083
rect 252 -1100 260 -1083
rect 294 -1100 302 -1083
rect 331 -1100 339 -1083
rect 373 -1100 381 -1083
rect -470 -1151 -453 -1120
rect 453 -1151 470 -1120
rect -470 -1168 -422 -1151
rect 422 -1168 470 -1151
<< viali >>
rect -372 1083 -338 1100
rect -293 1083 -259 1100
rect -214 1083 -180 1100
rect -135 1083 -101 1100
rect -56 1083 -22 1100
rect 23 1083 57 1100
rect 102 1083 136 1100
rect 181 1083 215 1100
rect 260 1083 294 1100
rect 339 1083 373 1100
rect -403 65 -386 1053
rect -324 65 -307 1053
rect -245 65 -228 1053
rect -166 65 -149 1053
rect -87 65 -70 1053
rect -8 65 9 1053
rect 71 65 88 1053
rect 150 65 167 1053
rect 229 65 246 1053
rect 308 65 325 1053
rect 387 65 404 1053
rect -372 18 -338 35
rect -293 18 -259 35
rect -214 18 -180 35
rect -135 18 -101 35
rect -56 18 -22 35
rect 23 18 57 35
rect 102 18 136 35
rect 181 18 215 35
rect 260 18 294 35
rect 339 18 373 35
rect -372 -35 -338 -18
rect -293 -35 -259 -18
rect -214 -35 -180 -18
rect -135 -35 -101 -18
rect -56 -35 -22 -18
rect 23 -35 57 -18
rect 102 -35 136 -18
rect 181 -35 215 -18
rect 260 -35 294 -18
rect 339 -35 373 -18
rect -403 -1053 -386 -65
rect -324 -1053 -307 -65
rect -245 -1053 -228 -65
rect -166 -1053 -149 -65
rect -87 -1053 -70 -65
rect -8 -1053 9 -65
rect 71 -1053 88 -65
rect 150 -1053 167 -65
rect 229 -1053 246 -65
rect 308 -1053 325 -65
rect 387 -1053 404 -65
rect -372 -1100 -338 -1083
rect -293 -1100 -259 -1083
rect -214 -1100 -180 -1083
rect -135 -1100 -101 -1083
rect -56 -1100 -22 -1083
rect 23 -1100 57 -1083
rect 102 -1100 136 -1083
rect 181 -1100 215 -1083
rect 260 -1100 294 -1083
rect 339 -1100 373 -1083
<< metal1 >>
rect -378 1100 -332 1103
rect -378 1083 -372 1100
rect -338 1083 -332 1100
rect -378 1080 -332 1083
rect -299 1100 -253 1103
rect -299 1083 -293 1100
rect -259 1083 -253 1100
rect -299 1080 -253 1083
rect -220 1100 -174 1103
rect -220 1083 -214 1100
rect -180 1083 -174 1100
rect -220 1080 -174 1083
rect -141 1100 -95 1103
rect -141 1083 -135 1100
rect -101 1083 -95 1100
rect -141 1080 -95 1083
rect -62 1100 -16 1103
rect -62 1083 -56 1100
rect -22 1083 -16 1100
rect -62 1080 -16 1083
rect 17 1100 63 1103
rect 17 1083 23 1100
rect 57 1083 63 1100
rect 17 1080 63 1083
rect 96 1100 142 1103
rect 96 1083 102 1100
rect 136 1083 142 1100
rect 96 1080 142 1083
rect 175 1100 221 1103
rect 175 1083 181 1100
rect 215 1083 221 1100
rect 175 1080 221 1083
rect 254 1100 300 1103
rect 254 1083 260 1100
rect 294 1083 300 1100
rect 254 1080 300 1083
rect 333 1100 379 1103
rect 333 1083 339 1100
rect 373 1083 379 1100
rect 333 1080 379 1083
rect -406 1053 -383 1059
rect -406 65 -403 1053
rect -386 65 -383 1053
rect -406 59 -383 65
rect -327 1053 -304 1059
rect -327 65 -324 1053
rect -307 65 -304 1053
rect -327 59 -304 65
rect -248 1053 -225 1059
rect -248 65 -245 1053
rect -228 65 -225 1053
rect -248 59 -225 65
rect -169 1053 -146 1059
rect -169 65 -166 1053
rect -149 65 -146 1053
rect -169 59 -146 65
rect -90 1053 -67 1059
rect -90 65 -87 1053
rect -70 65 -67 1053
rect -90 59 -67 65
rect -11 1053 13 1059
rect -11 65 -8 1053
rect 9 65 13 1053
rect -11 59 13 65
rect 68 1053 91 1059
rect 68 65 71 1053
rect 88 65 91 1053
rect 68 59 91 65
rect 147 1053 170 1059
rect 147 65 150 1053
rect 167 65 170 1053
rect 147 59 170 65
rect 226 1053 249 1059
rect 226 65 229 1053
rect 246 65 249 1053
rect 226 59 249 65
rect 305 1053 328 1059
rect 305 65 308 1053
rect 325 65 328 1053
rect 305 59 328 65
rect 384 1053 407 1059
rect 384 65 387 1053
rect 404 65 407 1053
rect 384 59 407 65
rect -378 35 -332 38
rect -378 18 -372 35
rect -338 18 -332 35
rect -378 15 -332 18
rect -299 35 -253 38
rect -299 18 -293 35
rect -259 18 -253 35
rect -299 15 -253 18
rect -220 35 -174 38
rect -220 18 -214 35
rect -180 18 -174 35
rect -220 15 -174 18
rect -141 35 -95 38
rect -141 18 -135 35
rect -101 18 -95 35
rect -141 15 -95 18
rect -62 35 -16 38
rect -62 18 -56 35
rect -22 18 -16 35
rect -62 15 -16 18
rect 17 35 63 38
rect 17 18 23 35
rect 57 18 63 35
rect 17 15 63 18
rect 96 35 142 38
rect 96 18 102 35
rect 136 18 142 35
rect 96 15 142 18
rect 175 35 221 38
rect 175 18 181 35
rect 215 18 221 35
rect 175 15 221 18
rect 254 35 300 38
rect 254 18 260 35
rect 294 18 300 35
rect 254 15 300 18
rect 333 35 379 38
rect 333 18 339 35
rect 373 18 379 35
rect 333 15 379 18
rect -378 -18 -332 -15
rect -378 -35 -372 -18
rect -338 -35 -332 -18
rect -378 -38 -332 -35
rect -299 -18 -253 -15
rect -299 -35 -293 -18
rect -259 -35 -253 -18
rect -299 -38 -253 -35
rect -220 -18 -174 -15
rect -220 -35 -214 -18
rect -180 -35 -174 -18
rect -220 -38 -174 -35
rect -141 -18 -95 -15
rect -141 -35 -135 -18
rect -101 -35 -95 -18
rect -141 -38 -95 -35
rect -62 -18 -16 -15
rect -62 -35 -56 -18
rect -22 -35 -16 -18
rect -62 -38 -16 -35
rect 17 -18 63 -15
rect 17 -35 23 -18
rect 57 -35 63 -18
rect 17 -38 63 -35
rect 96 -18 142 -15
rect 96 -35 102 -18
rect 136 -35 142 -18
rect 96 -38 142 -35
rect 175 -18 221 -15
rect 175 -35 181 -18
rect 215 -35 221 -18
rect 175 -38 221 -35
rect 254 -18 300 -15
rect 254 -35 260 -18
rect 294 -35 300 -18
rect 254 -38 300 -35
rect 333 -18 379 -15
rect 333 -35 339 -18
rect 373 -35 379 -18
rect 333 -38 379 -35
rect -406 -65 -383 -59
rect -406 -1053 -403 -65
rect -386 -1053 -383 -65
rect -406 -1059 -383 -1053
rect -327 -65 -304 -59
rect -327 -1053 -324 -65
rect -307 -1053 -304 -65
rect -327 -1059 -304 -1053
rect -248 -65 -225 -59
rect -248 -1053 -245 -65
rect -228 -1053 -225 -65
rect -248 -1059 -225 -1053
rect -169 -65 -146 -59
rect -169 -1053 -166 -65
rect -149 -1053 -146 -65
rect -169 -1059 -146 -1053
rect -90 -65 -67 -59
rect -90 -1053 -87 -65
rect -70 -1053 -67 -65
rect -90 -1059 -67 -1053
rect -11 -65 12 -59
rect -11 -1053 -8 -65
rect 9 -1053 12 -65
rect -11 -1059 12 -1053
rect 68 -65 91 -59
rect 68 -1053 71 -65
rect 88 -1053 91 -65
rect 68 -1059 91 -1053
rect 147 -65 170 -59
rect 147 -1053 150 -65
rect 167 -1053 170 -65
rect 147 -1059 170 -1053
rect 226 -65 249 -59
rect 226 -1053 229 -65
rect 246 -1053 249 -65
rect 226 -1059 249 -1053
rect 305 -65 328 -59
rect 305 -1053 308 -65
rect 325 -1053 328 -65
rect 305 -1059 328 -1053
rect 384 -65 407 -59
rect 384 -1053 387 -65
rect 404 -1053 407 -65
rect 384 -1059 407 -1053
rect -378 -1083 -332 -1080
rect -378 -1100 -372 -1083
rect -338 -1100 -332 -1083
rect -378 -1103 -332 -1100
rect -299 -1083 -253 -1080
rect -299 -1100 -293 -1083
rect -259 -1100 -253 -1083
rect -299 -1103 -253 -1100
rect -220 -1083 -174 -1080
rect -220 -1100 -214 -1083
rect -180 -1100 -174 -1083
rect -220 -1103 -174 -1100
rect -141 -1083 -95 -1080
rect -141 -1100 -135 -1083
rect -101 -1100 -95 -1083
rect -141 -1103 -95 -1100
rect -62 -1083 -16 -1080
rect -62 -1100 -56 -1083
rect -22 -1100 -16 -1083
rect -62 -1103 -16 -1100
rect 17 -1083 63 -1080
rect 17 -1100 23 -1083
rect 57 -1100 63 -1083
rect 17 -1103 63 -1100
rect 96 -1083 142 -1080
rect 96 -1100 102 -1083
rect 136 -1100 142 -1083
rect 96 -1103 142 -1100
rect 175 -1083 221 -1080
rect 175 -1100 181 -1083
rect 215 -1100 221 -1083
rect 175 -1103 221 -1100
rect 254 -1083 300 -1080
rect 254 -1100 260 -1083
rect 294 -1100 300 -1083
rect 254 -1103 300 -1100
rect 333 -1083 379 -1080
rect 333 -1100 339 -1083
rect 373 -1100 379 -1083
rect 333 -1103 379 -1100
<< properties >>
string FIXED_BBOX -462 -1160 462 1160
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.5 m 2 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
