magic
tech sky130A
timestamp 1644523392
<< nwell >>
rect -272 -648 272 648
<< mvpmos >>
rect -143 -500 -93 500
rect -64 -500 -14 500
rect 15 -500 65 500
rect 94 -500 144 500
<< mvpdiff >>
rect -172 494 -143 500
rect -172 -494 -166 494
rect -149 -494 -143 494
rect -172 -500 -143 -494
rect -93 494 -64 500
rect -93 -494 -87 494
rect -70 -494 -64 494
rect -93 -500 -64 -494
rect -14 494 15 500
rect -14 -494 -8 494
rect 9 -494 15 494
rect -14 -500 15 -494
rect 65 494 94 500
rect 65 -494 71 494
rect 88 -494 94 494
rect 65 -500 94 -494
rect 144 494 173 500
rect 144 -494 150 494
rect 167 -494 173 494
rect 144 -500 173 -494
<< mvpdiffc >>
rect -166 -494 -149 494
rect -87 -494 -70 494
rect -8 -494 9 494
rect 71 -494 88 494
rect 150 -494 167 494
<< mvnsubdiff >>
rect -239 609 239 615
rect -239 592 -185 609
rect 185 592 239 609
rect -239 586 239 592
rect -239 561 -210 586
rect -239 -561 -233 561
rect -216 -561 -210 561
rect 210 561 239 586
rect -239 -586 -210 -561
rect 210 -561 216 561
rect 233 -561 239 561
rect 210 -586 239 -561
rect -239 -592 239 -586
rect -239 -609 -185 -592
rect 185 -609 239 -592
rect -239 -615 239 -609
<< mvnsubdiffcont >>
rect -185 592 185 609
rect -233 -561 -216 561
rect 216 -561 233 561
rect -185 -609 185 -592
<< poly >>
rect -143 541 -93 549
rect -143 524 -135 541
rect -101 524 -93 541
rect -143 500 -93 524
rect -64 541 -14 549
rect -64 524 -56 541
rect -22 524 -14 541
rect -64 500 -14 524
rect 15 541 65 549
rect 15 524 23 541
rect 57 524 65 541
rect 15 500 65 524
rect 94 541 144 549
rect 94 524 102 541
rect 136 524 144 541
rect 94 500 144 524
rect -143 -524 -93 -500
rect -143 -541 -135 -524
rect -101 -541 -93 -524
rect -143 -549 -93 -541
rect -64 -524 -14 -500
rect -64 -541 -56 -524
rect -22 -541 -14 -524
rect -64 -549 -14 -541
rect 15 -524 65 -500
rect 15 -541 23 -524
rect 57 -541 65 -524
rect 15 -549 65 -541
rect 94 -524 144 -500
rect 94 -541 102 -524
rect 136 -541 144 -524
rect 94 -549 144 -541
<< polycont >>
rect -135 524 -101 541
rect -56 524 -22 541
rect 23 524 57 541
rect 102 524 136 541
rect -135 -541 -101 -524
rect -56 -541 -22 -524
rect 23 -541 57 -524
rect 102 -541 136 -524
<< locali >>
rect -233 592 -185 609
rect 185 592 233 609
rect -233 561 -216 592
rect 216 561 233 592
rect -143 524 -135 541
rect -101 524 -93 541
rect -64 524 -56 541
rect -22 524 -14 541
rect 15 524 23 541
rect 57 524 65 541
rect 94 524 102 541
rect 136 524 144 541
rect -166 494 -149 502
rect -166 -502 -149 -494
rect -87 494 -70 502
rect -87 -502 -70 -494
rect -8 494 9 502
rect -8 -502 9 -494
rect 71 494 88 502
rect 71 -502 88 -494
rect 150 494 167 502
rect 150 -502 167 -494
rect -143 -541 -135 -524
rect -101 -541 -93 -524
rect -64 -541 -56 -524
rect -22 -541 -14 -524
rect 15 -541 23 -524
rect 57 -541 65 -524
rect 94 -541 102 -524
rect 136 -541 144 -524
rect -233 -592 -216 -561
rect 216 -592 233 -561
rect -233 -609 -185 -592
rect 185 -609 233 -592
<< viali >>
rect -135 524 -101 541
rect -56 524 -22 541
rect 23 524 57 541
rect 102 524 136 541
rect -166 -494 -149 494
rect -87 -494 -70 494
rect -8 -494 9 494
rect 71 -494 88 494
rect 150 -494 167 494
rect -135 -541 -101 -524
rect -56 -541 -22 -524
rect 23 -541 57 -524
rect 102 -541 136 -524
<< metal1 >>
rect -141 541 -95 544
rect -141 524 -135 541
rect -101 524 -95 541
rect -141 521 -95 524
rect -62 541 -16 544
rect -62 524 -56 541
rect -22 524 -16 541
rect -62 521 -16 524
rect 17 541 63 544
rect 17 524 23 541
rect 57 524 63 541
rect 17 521 63 524
rect 96 541 142 544
rect 96 524 102 541
rect 136 524 142 541
rect 96 521 142 524
rect -169 494 -146 500
rect -169 -494 -166 494
rect -149 -494 -146 494
rect -169 -500 -146 -494
rect -90 494 -67 500
rect -90 -494 -87 494
rect -70 -494 -67 494
rect -90 -500 -67 -494
rect -11 494 12 500
rect -11 -494 -8 494
rect 9 -494 12 494
rect -11 -500 12 -494
rect 68 494 91 500
rect 68 -494 71 494
rect 88 -494 91 494
rect 68 -500 91 -494
rect 147 494 170 500
rect 147 -494 150 494
rect 167 -494 170 494
rect 147 -500 170 -494
rect -141 -524 -95 -521
rect -141 -541 -135 -524
rect -101 -541 -95 -524
rect -141 -544 -95 -541
rect -62 -524 -16 -521
rect -62 -541 -56 -524
rect -22 -541 -16 -524
rect -62 -544 -16 -541
rect 17 -524 63 -521
rect 17 -541 23 -524
rect 57 -541 63 -524
rect 17 -544 63 -541
rect 96 -524 142 -521
rect 96 -541 102 -524
rect 136 -541 142 -524
rect 96 -544 142 -541
<< properties >>
string FIXED_BBOX -225 -601 225 601
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
