magic
tech sky130A
magscale 1 2
timestamp 1721165872
<< nwell >>
rect -4532 -9608 -3054 -9512
rect -4558 -10622 -2972 -9608
rect -4364 -11930 -3372 -10622
rect -4490 -13308 -3188 -11930
rect -4330 -14242 -3338 -13308
rect -4330 -14362 -3848 -14242
rect -4330 -14618 -3864 -14362
<< locali >>
rect -3936 -9548 -3758 -9547
rect -3960 -9568 -3758 -9548
rect -1922 -9568 -1778 -9548
rect -5862 -9640 134 -9568
rect -5862 -11976 -5790 -9640
rect -3960 -11976 -3758 -9640
rect -5862 -12048 -3758 -11976
rect -5632 -12128 -3758 -12048
rect -5632 -13324 -5542 -12128
rect -4980 -13324 -4850 -12128
rect -5632 -13380 -4850 -13324
rect -5632 -13514 -4856 -13380
rect -5632 -14060 -5542 -13514
rect -4978 -14058 -4866 -13514
rect -3960 -14238 -3758 -12128
rect -1922 -11114 -1778 -9640
rect -1922 -11598 -1920 -11114
rect -1786 -11598 -1778 -11114
rect -1922 -13298 -1778 -11598
rect -1934 -13364 -1778 -13298
rect -1934 -13848 -1930 -13364
rect -1792 -13848 -1778 -13364
rect -1934 -13894 -1778 -13848
rect -1922 -14238 -1778 -13894
rect 62 -14238 134 -9640
rect -3960 -14310 134 -14238
rect -3960 -14410 128 -14310
rect -5590 -15278 -5500 -14656
rect -5068 -15178 -3766 -15094
rect -5078 -15212 -3766 -15178
rect -5078 -15278 -4952 -15212
rect -5590 -15284 -4952 -15278
rect -5590 -15396 -5392 -15284
rect -5130 -15322 -4952 -15284
rect -5130 -15396 -4954 -15322
rect -5590 -15408 -4954 -15396
rect -5590 -16582 -5500 -15408
rect -5070 -16582 -4954 -15408
rect -4064 -16558 -3766 -15212
rect -4064 -16582 122 -16558
rect -5590 -16702 122 -16582
rect -5510 -16706 122 -16702
rect -5263 -19058 -5161 -16706
rect -4110 -16759 122 -16706
rect -4110 -16772 -1778 -16759
rect -4110 -18054 -3768 -16772
rect -4066 -18420 -3768 -18054
rect -4118 -18620 -3768 -18420
rect -4110 -19058 -3768 -18620
rect -5263 -19078 -3768 -19058
rect -1920 -18156 -1778 -16772
rect -1920 -18640 -1918 -18156
rect -1786 -18640 -1778 -18156
rect -1920 -19078 -1778 -18640
rect 41 -19078 122 -16759
rect -5263 -19159 122 -19078
rect -5263 -19160 -4044 -19159
<< viali >>
rect -1920 -11598 -1786 -11114
rect -1930 -13848 -1792 -13364
rect -5392 -15396 -5130 -15284
rect -4118 -18420 -4066 -18054
rect -1918 -18640 -1786 -18156
<< metal1 >>
rect -5902 -9770 -4118 -9610
rect -3923 -9626 -3776 -9617
rect -5902 -11854 -5742 -9770
rect -5552 -10238 -5542 -9908
rect -5482 -10238 -5472 -9908
rect -5236 -10236 -5226 -9906
rect -5166 -10236 -5156 -9906
rect -4922 -10236 -4912 -9906
rect -4852 -10236 -4842 -9906
rect -4606 -10234 -4596 -9904
rect -4536 -10234 -4526 -9904
rect -4292 -10234 -4282 -9904
rect -4222 -10234 -4212 -9904
rect -3926 -9948 -3916 -9626
rect -3776 -9787 -91 -9633
rect -3776 -9948 -3766 -9787
rect -5712 -11678 -5702 -11348
rect -5642 -11678 -5632 -11348
rect -5396 -11676 -5386 -11346
rect -5326 -11676 -5316 -11346
rect -5082 -11678 -5072 -11348
rect -5012 -11678 -5002 -11348
rect -4762 -11680 -4752 -11350
rect -4692 -11680 -4682 -11350
rect -4446 -11680 -4436 -11350
rect -4376 -11680 -4366 -11350
rect -4130 -11680 -4120 -11350
rect -4060 -11680 -4050 -11350
rect -5902 -11962 -4100 -11854
rect -3923 -11874 -3769 -9948
rect -3554 -10772 -3544 -9902
rect -3418 -10772 -3408 -9902
rect -3236 -10772 -3226 -9902
rect -3100 -10772 -3090 -9902
rect -2922 -10774 -2912 -9904
rect -2786 -10774 -2776 -9904
rect -2606 -10774 -2596 -9904
rect -2470 -10774 -2460 -9904
rect -2288 -10774 -2278 -9904
rect -2152 -10774 -2142 -9904
rect -1550 -10772 -1544 -9902
rect -1418 -10772 -1412 -9902
rect -1232 -10772 -1226 -9902
rect -1100 -10772 -1094 -9902
rect -918 -10774 -912 -9904
rect -786 -10774 -780 -9904
rect -602 -10774 -596 -9904
rect -470 -10774 -464 -9904
rect -284 -10774 -278 -9904
rect -152 -10774 -146 -9904
rect -3708 -11760 -3698 -10890
rect -3572 -11760 -3562 -10890
rect -3390 -11760 -3380 -10890
rect -3254 -11760 -3244 -10890
rect -3076 -11762 -3066 -10892
rect -2940 -11762 -2930 -10892
rect -2760 -11762 -2750 -10892
rect -2624 -11762 -2614 -10892
rect -2442 -11762 -2432 -10892
rect -2306 -11762 -2296 -10892
rect -2128 -11762 -2118 -10892
rect -1992 -11762 -1982 -10892
rect -1926 -11114 -1778 -11102
rect -1930 -11598 -1920 -11114
rect -1786 -11598 -1778 -11114
rect -1926 -11610 -1778 -11598
rect -1704 -11760 -1698 -10890
rect -1572 -11760 -1566 -10890
rect -1386 -11760 -1380 -10890
rect -1254 -11760 -1248 -10890
rect -1072 -11762 -1066 -10892
rect -940 -11762 -934 -10892
rect -756 -11762 -750 -10892
rect -624 -11762 -618 -10892
rect -438 -11762 -432 -10892
rect -306 -11762 -300 -10892
rect -124 -11762 -118 -10892
rect 8 -11762 14 -10892
rect -5902 -14916 -5742 -11962
rect -3923 -12016 -87 -11874
rect -5906 -15120 -5896 -14916
rect -5756 -15120 -5742 -14916
rect -5902 -16668 -5742 -15120
rect -5612 -12282 -5132 -12230
rect -4718 -12278 -4106 -12228
rect -5612 -13166 -5560 -12282
rect -5458 -12680 -5448 -12450
rect -5388 -12680 -5378 -12450
rect -5146 -12680 -5136 -12450
rect -5076 -12680 -5066 -12450
rect -4764 -12672 -4754 -12442
rect -4694 -12672 -4684 -12442
rect -4446 -12678 -4436 -12448
rect -4376 -12678 -4366 -12448
rect -4134 -12678 -4124 -12448
rect -4064 -12678 -4054 -12448
rect -5302 -13056 -5292 -12926
rect -5232 -13056 -5222 -12926
rect -5612 -13218 -5122 -13166
rect -5612 -13536 -5560 -13218
rect -5612 -13588 -5082 -13536
rect -5612 -14964 -5560 -13588
rect -5450 -13670 -5398 -13588
rect -5464 -13800 -5454 -13670
rect -5394 -13800 -5384 -13670
rect -5302 -13798 -5292 -13668
rect -5232 -13798 -5222 -13668
rect -5134 -13672 -5082 -13588
rect -5146 -13802 -5136 -13672
rect -5076 -13802 -5066 -13672
rect -5328 -14860 -5220 -13880
rect -4604 -14248 -4594 -14018
rect -4534 -14248 -4524 -14018
rect -4284 -14246 -4274 -14016
rect -4214 -14246 -4204 -14016
rect -3923 -14108 -3769 -12016
rect -3554 -13008 -3544 -12138
rect -3418 -13008 -3408 -12138
rect -3236 -13008 -3226 -12138
rect -3100 -13008 -3090 -12138
rect -2922 -13010 -2912 -12140
rect -2786 -13010 -2776 -12140
rect -2606 -13010 -2596 -12140
rect -2470 -13010 -2460 -12140
rect -2288 -13010 -2278 -12140
rect -2152 -13010 -2142 -12140
rect -1550 -13008 -1544 -12138
rect -1418 -13008 -1412 -12138
rect -1232 -13008 -1226 -12138
rect -1100 -13008 -1094 -12138
rect -918 -13010 -912 -12140
rect -786 -13010 -780 -12140
rect -602 -13010 -596 -12140
rect -470 -13010 -464 -12140
rect -284 -13010 -278 -12140
rect -152 -13010 -146 -12140
rect -3708 -13996 -3698 -13126
rect -3572 -13996 -3562 -13126
rect -3390 -13996 -3380 -13126
rect -3254 -13996 -3244 -13126
rect -3076 -13998 -3066 -13128
rect -2940 -13998 -2930 -13128
rect -2760 -13998 -2750 -13128
rect -2624 -13998 -2614 -13128
rect -2442 -13998 -2432 -13128
rect -2306 -13998 -2296 -13128
rect -2128 -13998 -2118 -13128
rect -1992 -13998 -1982 -13128
rect -1936 -13364 -1786 -13352
rect -1940 -13848 -1930 -13364
rect -1792 -13848 -1786 -13364
rect -1936 -13860 -1786 -13848
rect -1704 -13996 -1698 -13126
rect -1572 -13996 -1566 -13126
rect -1386 -13996 -1380 -13126
rect -1254 -13996 -1248 -13126
rect -1072 -13998 -1066 -13128
rect -940 -13998 -934 -13128
rect -756 -13998 -750 -13128
rect -624 -13998 -618 -13128
rect -438 -13998 -432 -13128
rect -306 -13998 -300 -13128
rect -124 -13998 -118 -13128
rect 8 -13998 14 -13128
rect -3923 -14262 -91 -14108
rect -4692 -14418 -4118 -14362
rect -4616 -14520 -4526 -14418
rect -5056 -14540 -4526 -14520
rect -5056 -14662 -5046 -14540
rect -4938 -14662 -4526 -14540
rect -5056 -14678 -4526 -14662
rect -5612 -15016 -5348 -14964
rect -5216 -14968 -5114 -14894
rect -5612 -15506 -5560 -15016
rect -5178 -15236 -5114 -14968
rect -4616 -15135 -4526 -14678
rect -5400 -15248 -5114 -15236
rect -5400 -15284 -5388 -15248
rect -5400 -15396 -5392 -15284
rect -5400 -15402 -5388 -15396
rect -5126 -15402 -5114 -15248
rect -5400 -15420 -5114 -15402
rect -5059 -15225 -4526 -15135
rect -5612 -15558 -5236 -15506
rect -5612 -16420 -5560 -15558
rect -5059 -15853 -4969 -15225
rect -4616 -15304 -4526 -15225
rect -4794 -15360 -4220 -15304
rect -4704 -15724 -4694 -15494
rect -4634 -15724 -4624 -15494
rect -4386 -15724 -4376 -15494
rect -4316 -15724 -4306 -15494
rect -5205 -15943 -4969 -15853
rect -5410 -16318 -5400 -16084
rect -5330 -16318 -5320 -16084
rect -5612 -16472 -5226 -16420
rect -5031 -16424 -4981 -15943
rect -4860 -16316 -4850 -16086
rect -4790 -16316 -4780 -16086
rect -4540 -16314 -4530 -16084
rect -4470 -16314 -4460 -16084
rect -4230 -16320 -4220 -16090
rect -4160 -16320 -4150 -16090
rect -4078 -16320 -4068 -16090
rect -4008 -16320 -3998 -16090
rect -5031 -16474 -4210 -16424
rect -5902 -16802 -4124 -16668
rect -5902 -16858 -4122 -16802
rect -3923 -16806 -3769 -14262
rect -5298 -18924 -5190 -16858
rect -3923 -16888 -75 -16806
rect -3923 -16912 -3769 -16888
rect -4922 -17326 -4912 -16996
rect -4852 -17326 -4842 -16996
rect -4604 -17326 -4594 -16996
rect -4534 -17326 -4524 -16996
rect -4286 -17328 -4276 -16998
rect -4216 -17328 -4206 -16998
rect -3923 -17370 -3908 -16912
rect -3786 -17370 -3769 -16912
rect -4140 -18054 -4050 -18030
rect -4140 -18420 -4118 -18054
rect -4066 -18420 -4050 -18054
rect -4140 -18446 -4050 -18420
rect -5078 -18776 -5068 -18446
rect -5008 -18776 -4998 -18446
rect -4762 -18776 -4752 -18446
rect -4692 -18776 -4682 -18446
rect -4446 -18776 -4436 -18446
rect -4376 -18776 -4366 -18446
rect -4140 -18776 -4118 -18446
rect -4058 -18776 -4048 -18446
rect -4140 -18790 -4050 -18776
rect -5298 -19032 -4250 -18924
rect -3923 -18964 -3769 -17370
rect -3554 -17850 -3544 -16980
rect -3418 -17850 -3408 -16980
rect -3236 -17850 -3226 -16980
rect -3100 -17850 -3090 -16980
rect -2922 -17852 -2912 -16982
rect -2786 -17852 -2776 -16982
rect -2606 -17852 -2596 -16982
rect -2470 -17852 -2460 -16982
rect -2288 -17852 -2278 -16982
rect -2152 -17852 -2142 -16982
rect -1552 -17850 -1544 -16980
rect -1418 -17850 -1410 -16980
rect -1236 -17850 -1226 -16980
rect -1100 -17850 -1094 -16980
rect -920 -16982 -778 -16980
rect -920 -17852 -912 -16982
rect -786 -17850 -778 -16982
rect -604 -16982 -462 -16980
rect -786 -17852 -779 -17850
rect -604 -17852 -596 -16982
rect -470 -17850 -462 -16982
rect -288 -16982 -146 -16980
rect -470 -17852 -463 -17850
rect -288 -17852 -278 -16982
rect -152 -17852 -146 -16982
rect -3708 -18838 -3698 -17968
rect -3572 -18838 -3562 -17968
rect -3390 -18838 -3380 -17968
rect -3254 -18838 -3244 -17968
rect -3076 -18840 -3066 -17970
rect -2940 -18840 -2930 -17970
rect -2760 -18840 -2750 -17970
rect -2624 -18840 -2614 -17970
rect -2442 -18840 -2432 -17970
rect -2306 -18840 -2296 -17970
rect -2128 -18840 -2118 -17970
rect -1992 -18840 -1982 -17970
rect -1924 -18156 -1778 -18144
rect -1928 -18640 -1918 -18156
rect -1786 -18640 -1778 -18156
rect -1924 -18652 -1778 -18640
rect -1706 -18838 -1698 -17968
rect -1572 -18838 -1564 -17968
rect -1390 -18838 -1380 -17968
rect -1254 -18838 -1248 -17968
rect -1074 -17970 -932 -17968
rect -1074 -18840 -1066 -17970
rect -940 -18840 -932 -17970
rect -758 -17970 -616 -17968
rect -758 -18840 -750 -17970
rect -624 -18840 -616 -17970
rect -442 -17970 -300 -17968
rect -442 -18840 -432 -17970
rect -306 -18840 -300 -17970
rect -126 -17970 16 -17968
rect -126 -18840 -118 -17970
rect 8 -18840 16 -17970
rect -3923 -19118 -85 -18964
<< via1 >>
rect -5542 -10238 -5482 -9908
rect -5226 -10236 -5166 -9906
rect -4912 -10236 -4852 -9906
rect -4596 -10234 -4536 -9904
rect -4282 -10234 -4222 -9904
rect -3916 -9948 -3776 -9626
rect -5702 -11678 -5642 -11348
rect -5386 -11676 -5326 -11346
rect -5072 -11678 -5012 -11348
rect -4752 -11680 -4692 -11350
rect -4436 -11680 -4376 -11350
rect -4120 -11680 -4060 -11350
rect -3544 -10772 -3418 -9902
rect -3226 -10772 -3100 -9902
rect -2912 -10774 -2786 -9904
rect -2596 -10774 -2470 -9904
rect -2278 -10774 -2152 -9904
rect -1544 -10772 -1418 -9902
rect -1226 -10772 -1100 -9902
rect -912 -10774 -786 -9904
rect -596 -10774 -470 -9904
rect -278 -10774 -152 -9904
rect -3698 -11760 -3572 -10890
rect -3380 -11760 -3254 -10890
rect -3066 -11762 -2940 -10892
rect -2750 -11762 -2624 -10892
rect -2432 -11762 -2306 -10892
rect -2118 -11762 -1992 -10892
rect -1920 -11598 -1786 -11114
rect -1698 -11760 -1572 -10890
rect -1380 -11760 -1254 -10890
rect -1066 -11762 -940 -10892
rect -750 -11762 -624 -10892
rect -432 -11762 -306 -10892
rect -118 -11762 8 -10892
rect -5896 -15120 -5756 -14916
rect -5448 -12680 -5388 -12450
rect -5136 -12680 -5076 -12450
rect -4754 -12672 -4694 -12442
rect -4436 -12678 -4376 -12448
rect -4124 -12678 -4064 -12448
rect -5292 -13056 -5232 -12926
rect -5454 -13800 -5394 -13670
rect -5292 -13798 -5232 -13668
rect -5136 -13802 -5076 -13672
rect -4594 -14248 -4534 -14018
rect -4274 -14246 -4214 -14016
rect -3544 -13008 -3418 -12138
rect -3226 -13008 -3100 -12138
rect -2912 -13010 -2786 -12140
rect -2596 -13010 -2470 -12140
rect -2278 -13010 -2152 -12140
rect -1544 -13008 -1418 -12138
rect -1226 -13008 -1100 -12138
rect -912 -13010 -786 -12140
rect -596 -13010 -470 -12140
rect -278 -13010 -152 -12140
rect -3698 -13996 -3572 -13126
rect -3380 -13996 -3254 -13126
rect -3066 -13998 -2940 -13128
rect -2750 -13998 -2624 -13128
rect -2432 -13998 -2306 -13128
rect -2118 -13998 -1992 -13128
rect -1930 -13848 -1792 -13364
rect -1698 -13996 -1572 -13126
rect -1380 -13996 -1254 -13126
rect -1066 -13998 -940 -13128
rect -750 -13998 -624 -13128
rect -432 -13998 -306 -13128
rect -118 -13998 8 -13128
rect -5046 -14662 -4938 -14540
rect -5388 -15284 -5126 -15248
rect -5388 -15396 -5130 -15284
rect -5130 -15396 -5126 -15284
rect -5388 -15402 -5126 -15396
rect -4694 -15724 -4634 -15494
rect -4376 -15724 -4316 -15494
rect -5400 -16318 -5330 -16084
rect -4850 -16316 -4790 -16086
rect -4530 -16314 -4470 -16084
rect -4220 -16320 -4160 -16090
rect -4068 -16320 -4008 -16090
rect -4912 -17326 -4852 -16996
rect -4594 -17326 -4534 -16996
rect -4276 -17328 -4216 -16998
rect -3908 -17370 -3786 -16912
rect -5068 -18776 -5008 -18446
rect -4752 -18776 -4692 -18446
rect -4436 -18776 -4376 -18446
rect -4118 -18776 -4058 -18446
rect -3544 -17850 -3418 -16980
rect -3226 -17850 -3100 -16980
rect -2912 -17852 -2786 -16982
rect -2596 -17852 -2470 -16982
rect -2278 -17852 -2152 -16982
rect -1544 -17850 -1418 -16980
rect -1226 -17850 -1100 -16980
rect -912 -17852 -786 -16982
rect -596 -17852 -470 -16982
rect -278 -17852 -152 -16982
rect -3698 -18838 -3572 -17968
rect -3380 -18838 -3254 -17968
rect -3066 -18840 -2940 -17970
rect -2750 -18840 -2624 -17970
rect -2432 -18840 -2306 -17970
rect -2118 -18840 -1992 -17970
rect -1900 -18638 -1786 -18176
rect -1698 -18838 -1572 -17968
rect -1380 -18838 -1254 -17968
rect -1066 -18840 -940 -17970
rect -750 -18840 -624 -17970
rect -432 -18840 -306 -17970
rect -118 -18840 8 -17970
<< metal2 >>
rect -3932 -9616 -3848 -9612
rect -3932 -9626 -3776 -9616
rect -5542 -9908 -5482 -9898
rect -5226 -9906 -5166 -9896
rect -5482 -10208 -5226 -9924
rect -5542 -10248 -5482 -10238
rect -4912 -9906 -4852 -9896
rect -5166 -10208 -4912 -9924
rect -5226 -10246 -5166 -10236
rect -4596 -9904 -4536 -9894
rect -4852 -10208 -4596 -9924
rect -4912 -10246 -4852 -10236
rect -4282 -9904 -4222 -9894
rect -4536 -10208 -4282 -9924
rect -4596 -10244 -4536 -10234
rect -3932 -9924 -3916 -9626
rect -4222 -9948 -3916 -9924
rect -4222 -10208 -3776 -9948
rect -3544 -9902 -3418 -9892
rect -4282 -10244 -4222 -10234
rect -3226 -9902 -3100 -9892
rect -3418 -10614 -3226 -10080
rect -3544 -10782 -3418 -10772
rect -2912 -9904 -2786 -9894
rect -3100 -10614 -2912 -10080
rect -3226 -10782 -3100 -10772
rect -2596 -9904 -2470 -9894
rect -2786 -10614 -2596 -10080
rect -2912 -10784 -2786 -10774
rect -2278 -9904 -2152 -9894
rect -2470 -10614 -2278 -10080
rect -2596 -10784 -2470 -10774
rect -1544 -9902 -1418 -9892
rect -2152 -10092 -1544 -10080
rect -1226 -9902 -1100 -9892
rect -1418 -10092 -1226 -10080
rect -912 -9904 -786 -9894
rect -1100 -10092 -912 -10080
rect -596 -9904 -470 -9894
rect -786 -10092 -596 -10080
rect -278 -9904 -152 -9894
rect -470 -10092 -278 -10080
rect -2152 -10602 -1590 -10092
rect -2152 -10614 -1544 -10602
rect -2278 -10784 -2152 -10774
rect -1418 -10614 -1226 -10602
rect -1544 -10782 -1418 -10772
rect -1100 -10614 -912 -10602
rect -1226 -10782 -1100 -10772
rect -786 -10614 -596 -10602
rect -912 -10784 -786 -10774
rect -470 -10614 -278 -10602
rect -596 -10784 -470 -10774
rect -152 -10614 -134 -10080
rect -278 -10784 -152 -10774
rect -3890 -10890 -3730 -10888
rect -3698 -10890 -3572 -10880
rect -5702 -11348 -5642 -11338
rect -5386 -11346 -5326 -11336
rect -5642 -11656 -5386 -11372
rect -5702 -11688 -5642 -11678
rect -5072 -11348 -5012 -11338
rect -5326 -11656 -5072 -11372
rect -5386 -11686 -5326 -11676
rect -4752 -11350 -4692 -11340
rect -5012 -11656 -4752 -11372
rect -5072 -11688 -5012 -11678
rect -4436 -11350 -4376 -11340
rect -4692 -11656 -4436 -11372
rect -4752 -11690 -4692 -11680
rect -4120 -11350 -4060 -11340
rect -4376 -11656 -4120 -11372
rect -4436 -11690 -4376 -11680
rect -3890 -11372 -3698 -10890
rect -3380 -10890 -3254 -10880
rect -3572 -11234 -3380 -11114
rect -3066 -10892 -2940 -10882
rect -3254 -11234 -3066 -11114
rect -2750 -10892 -2624 -10882
rect -2940 -11234 -2750 -11114
rect -2432 -10892 -2306 -10882
rect -2624 -11234 -2432 -11114
rect -2118 -10892 -1992 -10882
rect -1698 -10890 -1572 -10880
rect -2306 -11234 -2118 -11114
rect -1920 -11114 -1782 -11104
rect -1736 -11114 -1698 -10890
rect -1992 -11234 -1920 -11114
rect -4060 -11656 -3698 -11372
rect -4120 -11690 -4060 -11680
rect -3889 -11760 -3698 -11656
rect -3572 -11600 -3380 -11548
rect -3889 -11770 -3572 -11760
rect -3254 -11600 -3066 -11548
rect -3380 -11770 -3254 -11760
rect -2940 -11600 -2750 -11548
rect -3889 -11772 -3654 -11770
rect -3066 -11772 -2940 -11762
rect -2624 -11600 -2432 -11548
rect -2750 -11772 -2624 -11762
rect -2306 -11600 -2118 -11548
rect -2432 -11772 -2306 -11762
rect -1992 -11598 -1920 -11548
rect -1786 -11598 -1698 -11114
rect -1992 -11600 -1698 -11598
rect -1920 -11608 -1782 -11600
rect -2118 -11772 -1992 -11762
rect -1736 -11760 -1698 -11600
rect -1380 -10890 -1254 -10880
rect -1572 -11600 -1380 -11114
rect -1736 -11770 -1572 -11760
rect -1066 -10892 -940 -10882
rect -1254 -11600 -1066 -11114
rect -1380 -11770 -1254 -11760
rect -750 -10892 -624 -10882
rect -940 -11600 -750 -11114
rect -1736 -11772 -1654 -11770
rect -1066 -11772 -940 -11762
rect -432 -10892 -306 -10882
rect -624 -11600 -432 -11114
rect -750 -11772 -624 -11762
rect -118 -10892 8 -10882
rect -306 -11600 -118 -11114
rect -432 -11772 -306 -11762
rect 8 -11600 28 -11114
rect -118 -11772 8 -11762
rect -5448 -12450 -5388 -12440
rect -5136 -12450 -5076 -12440
rect -5388 -12650 -5136 -12472
rect -5448 -12690 -5388 -12680
rect -4754 -12442 -4694 -12432
rect -5076 -12650 -4754 -12472
rect -5136 -12690 -5076 -12680
rect -5292 -12926 -5232 -12916
rect -5606 -13036 -5292 -12958
rect -5606 -14563 -5528 -13036
rect -5292 -13066 -5232 -13056
rect -4977 -13403 -4899 -12650
rect -4436 -12448 -4376 -12438
rect -4694 -12650 -4436 -12472
rect -4754 -12682 -4694 -12672
rect -4124 -12448 -4064 -12438
rect -4376 -12650 -4124 -12472
rect -4436 -12688 -4376 -12678
rect -3889 -12472 -3811 -11772
rect -4064 -12650 -3811 -12472
rect -3544 -12138 -3418 -12128
rect -4124 -12688 -4064 -12678
rect -3226 -12138 -3100 -12128
rect -3418 -12806 -3226 -12272
rect -3544 -13018 -3418 -13008
rect -2912 -12140 -2786 -12130
rect -3100 -12806 -2912 -12272
rect -3226 -13018 -3100 -13008
rect -2596 -12140 -2470 -12130
rect -2786 -12806 -2596 -12272
rect -2912 -13020 -2786 -13010
rect -2278 -12140 -2152 -12130
rect -2470 -12806 -2278 -12272
rect -2596 -13020 -2470 -13010
rect -1544 -12138 -1418 -12128
rect -2152 -12284 -1544 -12272
rect -1226 -12138 -1100 -12128
rect -1418 -12284 -1226 -12272
rect -912 -12140 -786 -12130
rect -1100 -12284 -912 -12272
rect -596 -12140 -470 -12130
rect -786 -12284 -596 -12272
rect -278 -12140 -152 -12130
rect -470 -12284 -278 -12272
rect -2152 -12794 -1590 -12284
rect -2152 -12806 -1544 -12794
rect -2278 -13020 -2152 -13010
rect -1418 -12806 -1226 -12794
rect -1544 -13018 -1418 -13008
rect -1100 -12806 -912 -12794
rect -1226 -13018 -1100 -13008
rect -786 -12806 -596 -12794
rect -912 -13020 -786 -13010
rect -470 -12806 -278 -12794
rect -596 -13020 -470 -13010
rect -152 -12806 -124 -12272
rect -278 -13020 -152 -13010
rect -5303 -13481 -4899 -13403
rect -3698 -13126 -3572 -13116
rect -5454 -13670 -5394 -13660
rect -5454 -13810 -5394 -13800
rect -5303 -13668 -5225 -13481
rect -3380 -13126 -3254 -13116
rect -3572 -13488 -3380 -13366
rect -3066 -13128 -2940 -13118
rect -3254 -13488 -3066 -13366
rect -2750 -13128 -2624 -13118
rect -2940 -13488 -2750 -13366
rect -2432 -13128 -2306 -13118
rect -2624 -13488 -2432 -13366
rect -2118 -13128 -1992 -13118
rect -2306 -13488 -2118 -13366
rect -1698 -13126 -1572 -13116
rect -1930 -13364 -1792 -13354
rect -1992 -13488 -1930 -13366
rect -5303 -13798 -5292 -13668
rect -5232 -13798 -5225 -13668
rect -5303 -13815 -5225 -13798
rect -5136 -13672 -5076 -13662
rect -5136 -13812 -5076 -13802
rect -3572 -13852 -3380 -13802
rect -3698 -14006 -3572 -13996
rect -3254 -13852 -3066 -13802
rect -3380 -14006 -3254 -13996
rect -2940 -13852 -2750 -13802
rect -4594 -14018 -4534 -14008
rect -4274 -14016 -4214 -14006
rect -3066 -14008 -2940 -13998
rect -2624 -13852 -2432 -13802
rect -2750 -14008 -2624 -13998
rect -2306 -13852 -2118 -13802
rect -2432 -14008 -2306 -13998
rect -1992 -13848 -1930 -13802
rect -1792 -13848 -1698 -13366
rect -1992 -13852 -1698 -13848
rect -1930 -13858 -1792 -13852
rect -2118 -14008 -1992 -13998
rect -1380 -13126 -1254 -13116
rect -1572 -13852 -1380 -13366
rect -1698 -14006 -1572 -13996
rect -1066 -13128 -940 -13118
rect -1254 -13852 -1066 -13366
rect -1380 -14006 -1254 -13996
rect -750 -13128 -624 -13118
rect -940 -13852 -750 -13366
rect -1066 -14008 -940 -13998
rect -432 -13128 -306 -13118
rect -624 -13852 -432 -13366
rect -750 -14008 -624 -13998
rect -118 -13128 8 -13118
rect -306 -13852 -118 -13366
rect -432 -14008 -306 -13998
rect 8 -13852 28 -13366
rect -118 -14008 8 -13998
rect -4534 -14228 -4274 -14034
rect -4594 -14258 -4534 -14248
rect -5046 -14540 -4938 -14530
rect -5606 -14641 -5046 -14563
rect -5046 -14672 -4938 -14662
rect -5896 -14916 -5756 -14906
rect -4479 -14979 -4393 -14228
rect -4274 -14256 -4214 -14246
rect -5756 -15065 -4393 -14979
rect -5896 -15130 -5756 -15120
rect -5400 -15248 -5114 -15236
rect -5400 -15402 -5388 -15248
rect -5126 -15402 -5114 -15248
rect -5400 -15420 -5114 -15402
rect -5398 -16074 -5336 -15420
rect -4479 -15484 -4393 -15065
rect -4694 -15494 -4634 -15484
rect -4479 -15494 -4316 -15484
rect -4479 -15514 -4376 -15494
rect -4634 -15700 -4376 -15514
rect -4694 -15734 -4634 -15724
rect -4376 -15734 -4316 -15724
rect -5400 -16084 -5330 -16074
rect -5414 -16296 -5400 -16110
rect -4850 -16086 -4790 -16076
rect -5330 -16296 -4850 -16110
rect -5400 -16328 -5330 -16318
rect -5089 -18166 -5003 -16296
rect -4530 -16084 -4470 -16074
rect -4790 -16296 -4530 -16110
rect -4850 -16326 -4790 -16316
rect -4220 -16090 -4160 -16080
rect -4470 -16296 -4220 -16110
rect -4530 -16324 -4470 -16314
rect -4068 -16090 -4008 -16080
rect -4084 -16114 -4068 -16110
rect -4101 -16115 -4068 -16114
rect -4160 -16289 -4068 -16115
rect -4084 -16296 -4068 -16289
rect -4220 -16330 -4160 -16320
rect -4008 -16289 -3992 -16115
rect -4068 -16330 -4008 -16320
rect -3908 -16912 -3786 -16902
rect -4912 -16996 -4852 -16986
rect -4932 -17312 -4912 -17006
rect -4594 -16996 -4534 -16986
rect -4852 -17312 -4594 -17006
rect -4912 -17336 -4852 -17326
rect -4276 -16998 -4216 -16988
rect -4534 -17312 -4276 -17006
rect -4594 -17336 -4534 -17326
rect -4216 -17312 -3908 -17006
rect -4276 -17338 -4216 -17328
rect -3908 -17380 -3786 -17370
rect -3544 -16980 -3418 -16970
rect -3226 -16980 -3100 -16970
rect -3418 -17668 -3226 -17134
rect -3544 -17860 -3418 -17850
rect -2912 -16982 -2786 -16972
rect -3100 -17668 -2912 -17134
rect -3226 -17860 -3100 -17850
rect -2596 -16982 -2470 -16972
rect -2786 -17668 -2596 -17134
rect -2912 -17862 -2786 -17852
rect -2278 -16982 -2152 -16972
rect -2470 -17668 -2278 -17134
rect -2596 -17862 -2470 -17852
rect -1544 -16980 -1418 -16970
rect -2152 -17140 -1544 -17134
rect -1226 -16980 -1100 -16970
rect -1418 -17140 -1226 -17134
rect -912 -16982 -786 -16972
rect -1100 -17140 -912 -17134
rect -596 -16982 -470 -16972
rect -786 -17140 -596 -17134
rect -278 -16982 -152 -16972
rect -470 -17140 -278 -17134
rect -2152 -17650 -1588 -17140
rect -2152 -17668 -1544 -17650
rect -2278 -17862 -2152 -17852
rect -1418 -17668 -1226 -17650
rect -1544 -17860 -1418 -17850
rect -1100 -17668 -912 -17650
rect -1226 -17860 -1100 -17850
rect -786 -17668 -596 -17650
rect -912 -17862 -786 -17852
rect -470 -17668 -278 -17650
rect -596 -17862 -470 -17852
rect -152 -17668 -118 -17134
rect -278 -17862 -152 -17852
rect -3698 -17968 -3572 -17958
rect -5089 -18320 -3698 -18166
rect -3380 -17968 -3254 -17958
rect -3572 -18320 -3380 -18166
rect -3066 -17970 -2940 -17960
rect -5089 -18446 -5050 -18320
rect -5089 -18470 -5068 -18446
rect -5092 -18762 -5068 -18470
rect -5089 -18776 -5068 -18762
rect -5008 -18762 -4752 -18634
rect -5008 -18776 -5003 -18762
rect -5089 -18781 -5003 -18776
rect -4692 -18762 -4436 -18634
rect -5068 -18786 -5008 -18781
rect -4752 -18786 -4692 -18776
rect -4376 -18762 -4118 -18634
rect -4436 -18786 -4376 -18776
rect -4058 -18762 -3698 -18634
rect -4118 -18786 -4058 -18776
rect -3572 -18652 -3380 -18634
rect -3698 -18848 -3572 -18838
rect -3254 -18652 -3066 -18166
rect -3380 -18848 -3254 -18838
rect -2750 -17970 -2624 -17960
rect -2940 -18652 -2750 -18166
rect -3066 -18850 -2940 -18840
rect -2432 -17970 -2306 -17960
rect -2624 -18652 -2432 -18166
rect -2750 -18850 -2624 -18840
rect -2118 -17970 -1992 -17960
rect -2306 -18652 -2118 -18166
rect -2432 -18850 -2306 -18840
rect -1698 -17968 -1572 -17958
rect -1992 -18176 -1698 -18166
rect -1992 -18638 -1900 -18176
rect -1786 -18638 -1698 -18176
rect -1992 -18652 -1698 -18638
rect -2118 -18850 -1992 -18840
rect -1380 -17968 -1254 -17958
rect -1572 -18652 -1380 -18166
rect -1698 -18848 -1572 -18838
rect -1066 -17970 -940 -17960
rect -1254 -18652 -1066 -18166
rect -1380 -18848 -1254 -18838
rect -750 -17970 -624 -17960
rect -940 -18652 -750 -18166
rect -1066 -18850 -940 -18840
rect -432 -17970 -306 -17960
rect -624 -18652 -432 -18166
rect -750 -18850 -624 -18840
rect -118 -17970 8 -17960
rect -306 -18652 -118 -18166
rect -432 -18850 -306 -18840
rect 8 -18652 40 -18166
rect -118 -18850 8 -18840
<< via2 >>
rect -1590 -10602 -1544 -10092
rect -1544 -10602 -1418 -10092
rect -1418 -10602 -1226 -10092
rect -1226 -10602 -1100 -10092
rect -1100 -10602 -912 -10092
rect -912 -10602 -786 -10092
rect -786 -10602 -596 -10092
rect -596 -10602 -470 -10092
rect -470 -10602 -278 -10092
rect -278 -10602 -168 -10092
rect -3614 -11548 -3572 -11234
rect -3572 -11548 -3380 -11234
rect -3380 -11548 -3254 -11234
rect -3254 -11548 -3066 -11234
rect -3066 -11548 -2940 -11234
rect -2940 -11548 -2750 -11234
rect -2750 -11548 -2624 -11234
rect -2624 -11548 -2432 -11234
rect -2432 -11548 -2306 -11234
rect -2306 -11548 -2118 -11234
rect -2118 -11548 -1992 -11234
rect -1992 -11548 -1920 -11234
rect -1920 -11548 -1896 -11234
rect -1590 -12794 -1544 -12284
rect -1544 -12794 -1418 -12284
rect -1418 -12794 -1226 -12284
rect -1226 -12794 -1100 -12284
rect -1100 -12794 -912 -12284
rect -912 -12794 -786 -12284
rect -786 -12794 -596 -12284
rect -596 -12794 -470 -12284
rect -470 -12794 -278 -12284
rect -278 -12794 -168 -12284
rect -3608 -13802 -3572 -13488
rect -3572 -13802 -3380 -13488
rect -3380 -13802 -3254 -13488
rect -3254 -13802 -3066 -13488
rect -3066 -13802 -2940 -13488
rect -2940 -13802 -2750 -13488
rect -2750 -13802 -2624 -13488
rect -2624 -13802 -2432 -13488
rect -2432 -13802 -2306 -13488
rect -2306 -13802 -2118 -13488
rect -2118 -13802 -1992 -13488
rect -1992 -13802 -1930 -13488
rect -1930 -13802 -1914 -13488
rect -1588 -17650 -1544 -17140
rect -1544 -17650 -1418 -17140
rect -1418 -17650 -1226 -17140
rect -1226 -17650 -1100 -17140
rect -1100 -17650 -912 -17140
rect -912 -17650 -786 -17140
rect -786 -17650 -596 -17140
rect -596 -17650 -470 -17140
rect -470 -17650 -278 -17140
rect -278 -17650 -166 -17140
rect -5050 -18446 -3698 -18320
rect -5050 -18634 -5008 -18446
rect -5008 -18634 -4752 -18446
rect -4752 -18634 -4692 -18446
rect -4692 -18634 -4436 -18446
rect -4436 -18634 -4376 -18446
rect -4376 -18634 -4118 -18446
rect -4118 -18634 -4058 -18446
rect -4058 -18634 -3698 -18446
rect -3698 -18634 -3572 -18320
rect -3572 -18634 -3380 -18320
rect -3380 -18634 -3292 -18320
<< metal3 >>
rect -3644 -11234 -1880 -8966
rect -1594 -10087 -156 -8926
rect -1600 -10092 -156 -10087
rect -1600 -10602 -1590 -10092
rect -168 -10602 -156 -10092
rect -1600 -10607 -156 -10602
rect -3644 -11548 -3614 -11234
rect -1896 -11548 -1880 -11234
rect -3644 -13488 -1880 -11548
rect -1594 -12279 -156 -10607
rect -1600 -12284 -156 -12279
rect -1600 -12794 -1590 -12284
rect -168 -12794 -156 -12284
rect -1600 -12799 -156 -12794
rect -3644 -13802 -3608 -13488
rect -1914 -13802 -1880 -13488
rect -3644 -14242 -1880 -13802
rect -5056 -18320 -3278 -18310
rect -5056 -18634 -5050 -18320
rect -3292 -18634 -3278 -18320
rect -5056 -18640 -3278 -18634
rect -5050 -19824 -3278 -18640
rect -3154 -19828 -1880 -14242
rect -1594 -14545 -156 -12799
rect -1594 -15065 -152 -14545
rect -1594 -17135 -156 -15065
rect -1598 -17140 -156 -17135
rect -1598 -17650 -1588 -17140
rect -166 -17650 -156 -17140
rect -1598 -17655 -156 -17650
rect -1594 -19824 -156 -17655
use sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3  sky130_fd_pr__nfet_g5v0d10v5_MJGQJ3_0 paramcells
timestamp 1644523392
transform 1 0 -5280 0 1 -15988
box -278 -658 278 658
use sky130_fd_pr__nfet_g5v0d10v5_QABAEG  sky130_fd_pr__nfet_g5v0d10v5_QABAEG_0 paramcells
timestamp 1644523392
transform 1 0 -4505 0 1 -15888
box -514 -758 514 758
use sky130_fd_pr__nfet_g5v0d10v5_QCNVDG  sky130_fd_pr__nfet_g5v0d10v5_QCNVDG_0 paramcells
timestamp 1721163516
transform 1 0 -4640 0 1 -17889
box -594 -1258 594 1258
use sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ  sky130_fd_pr__nfet_g5v0d10v5_RX3AJQ_0 paramcells
timestamp 1644523392
transform 1 0 -5280 0 1 -14990
box -278 -358 278 358
use sky130_fd_pr__nfet_g5v0d10v5_YSH3F7  sky130_fd_pr__nfet_g5v0d10v5_YSH3F7_0 paramcells
timestamp 1721163516
transform 1 0 -843 0 1 -17928
box -989 -1258 989 1258
use sky130_fd_pr__nfet_g5v0d10v5_YSH3F7  sky130_fd_pr__nfet_g5v0d10v5_YSH3F7_1
timestamp 1721163516
transform 1 0 -2843 0 1 -17928
box -989 -1258 989 1258
use sky130_fd_pr__pfet_g5v0d10v5_3QQKN5  sky130_fd_pr__pfet_g5v0d10v5_3QQKN5_1 paramcells
timestamp 1644523392
transform 1 0 -5262 0 1 -12726
box -386 -696 386 696
use sky130_fd_pr__pfet_g5v0d10v5_54K6JW  sky130_fd_pr__pfet_g5v0d10v5_54K6JW_0 paramcells
timestamp 1721163516
transform 1 0 -2843 0 1 -11947
box -1019 -2415 1019 2415
use sky130_fd_pr__pfet_g5v0d10v5_54K6JW  sky130_fd_pr__pfet_g5v0d10v5_54K6JW_1
timestamp 1721163516
transform 1 0 -843 0 1 -11947
box -1019 -2415 1019 2415
use sky130_fd_pr__pfet_g5v0d10v5_CYU746  sky130_fd_pr__pfet_g5v0d10v5_CYU746_0 paramcells
timestamp 1721163516
transform 1 0 -4881 0 1 -10809
box -1019 -1297 1019 1297
use sky130_fd_pr__pfet_g5v0d10v5_HKUKAU  sky130_fd_pr__pfet_g5v0d10v5_HKUKAU_0 paramcells
timestamp 1644523392
transform 1 0 -5263 0 1 -13774
box -386 -362 386 362
use sky130_fd_pr__pfet_g5v0d10v5_WECJAU  sky130_fd_pr__pfet_g5v0d10v5_WECJAU_0 paramcells
timestamp 1644523392
transform 1 0 -4407 0 1 -13325
box -544 -1296 544 1296
<< labels >>
rlabel metal1 -5328 -14860 -5220 -13880 1 in
port 1 n
rlabel metal1 -5612 -15558 -5560 -13166 1 drv1
rlabel metal2 -5606 -14641 -4938 -14563 1 drv2
rlabel metal1 -5902 -16858 -5742 -15120 1 crosscon
port 2 n
rlabel metal1 -3923 -16912 -3769 -9948 1 drv4
rlabel metal3 -3644 -14242 -2400 -13802 1 vdd_hi
port 4 n
rlabel metal3 -1594 -14550 -676 -12794 1 out
port 3 n
rlabel metal3 -4974 -19824 -3724 -18634 1 vss
port 5 n
<< end >>
