magic
tech sky130A
timestamp 1644523392
<< nwell >>
rect -193 -181 193 181
<< mvpmos >>
rect -64 -32 -14 68
rect 15 -32 65 68
<< mvpdiff >>
rect -93 62 -64 68
rect -93 -26 -87 62
rect -70 -26 -64 62
rect -93 -32 -64 -26
rect -14 62 15 68
rect -14 -26 -8 62
rect 9 -26 15 62
rect -14 -32 15 -26
rect 65 62 94 68
rect 65 -26 71 62
rect 88 -26 94 62
rect 65 -32 94 -26
<< mvpdiffc >>
rect -87 -26 -70 62
rect -8 -26 9 62
rect 71 -26 88 62
<< mvnsubdiff >>
rect -160 142 160 148
rect -160 125 -106 142
rect 106 125 160 142
rect -160 119 160 125
rect -160 94 -131 119
rect -160 -94 -154 94
rect -137 -94 -131 94
rect 131 94 160 119
rect -160 -119 -131 -94
rect 131 -94 137 94
rect 154 -94 160 94
rect 131 -119 160 -94
rect -160 -125 160 -119
rect -160 -142 -106 -125
rect 106 -142 160 -125
rect -160 -148 160 -142
<< mvnsubdiffcont >>
rect -106 125 106 142
rect -154 -94 -137 94
rect 137 -94 154 94
rect -106 -142 106 -125
<< poly >>
rect -64 68 -14 81
rect 15 68 65 81
rect -64 -56 -14 -32
rect -64 -73 -56 -56
rect -22 -73 -14 -56
rect -64 -81 -14 -73
rect 15 -56 65 -32
rect 15 -73 23 -56
rect 57 -73 65 -56
rect 15 -81 65 -73
<< polycont >>
rect -56 -73 -22 -56
rect 23 -73 57 -56
<< locali >>
rect -154 125 -106 142
rect 106 125 154 142
rect -154 94 -137 125
rect 137 94 154 125
rect -87 62 -70 70
rect -87 -34 -70 -26
rect -8 62 9 70
rect -8 -34 9 -26
rect 71 62 88 70
rect 71 -34 88 -26
rect -64 -73 -56 -56
rect -22 -73 -14 -56
rect 15 -73 23 -56
rect 57 -73 65 -56
rect -154 -125 -137 -94
rect 137 -125 154 -94
rect -154 -142 -106 -125
rect 106 -142 154 -125
<< viali >>
rect -87 -26 -70 62
rect -8 -26 9 62
rect 71 -26 88 62
rect -56 -73 -22 -56
rect 23 -73 57 -56
<< metal1 >>
rect -90 62 -67 68
rect -90 -26 -87 62
rect -70 -26 -67 62
rect -90 -32 -67 -26
rect -11 62 12 68
rect -11 -26 -8 62
rect 9 -26 12 62
rect -11 -32 12 -26
rect 68 62 91 68
rect 68 -26 71 62
rect 88 -26 91 62
rect 68 -32 91 -26
rect -62 -56 -16 -53
rect -62 -73 -56 -56
rect -22 -73 -16 -56
rect -62 -76 -16 -73
rect 17 -56 63 -53
rect 17 -73 23 -56
rect 57 -73 63 -56
rect 17 -76 63 -73
<< properties >>
string FIXED_BBOX -146 -133 146 133
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
