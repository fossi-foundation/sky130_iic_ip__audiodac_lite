magic
tech sky130A
magscale 1 2
timestamp 1747753545
<< dnwell >>
rect -206 -190 9522 28568
<< nwell >>
rect -316 28362 9632 28678
rect -316 16792 47 28362
rect 2533 28114 2853 28362
rect 2521 28094 2853 28114
rect 2521 27358 2811 28094
rect 2541 26124 2809 27358
rect 2541 24140 2807 26124
rect 2527 23558 2849 24140
rect 2527 23536 3061 23558
rect 2551 23530 3061 23536
rect -316 11594 0 16792
rect -316 16 27 11594
rect 2529 4836 2621 4838
rect 2529 4818 3047 4836
rect 2529 4808 2833 4818
rect 2495 1242 2833 4808
rect 2501 218 2833 1242
rect 2501 46 2897 218
rect 2435 16 2969 46
rect 9316 16 9632 28362
rect -316 -300 9632 16
<< mvnsubdiff >>
rect -249 28591 9565 28611
rect -249 28557 -169 28591
rect 9485 28557 9565 28591
rect -249 28537 9565 28557
rect -249 28531 -175 28537
rect -249 -153 -229 28531
rect -195 -153 -175 28531
rect -249 -159 -175 -153
rect 9491 28531 9565 28537
rect 9491 -153 9511 28531
rect 9545 -153 9565 28531
rect 9491 -159 9565 -153
rect -249 -179 9565 -159
rect -249 -213 -169 -179
rect 9485 -213 9565 -179
rect -249 -233 9565 -213
<< mvnsubdiffcont >>
rect -169 28557 9485 28591
rect -229 -153 -195 28531
rect 9511 -153 9545 28531
rect -169 -213 9485 -179
<< locali >>
rect -249 28602 9567 28621
rect -249 28591 -148 28602
rect 9456 28591 9567 28602
rect -249 28557 -169 28591
rect 9485 28557 9567 28591
rect -249 28550 -148 28557
rect 9456 28550 9567 28557
rect -249 28531 9567 28550
rect -249 28494 -229 28531
rect -195 28503 9511 28531
rect -195 28494 -131 28503
rect -249 -86 -238 28494
rect -186 -86 -131 28494
rect 96 28340 184 28503
rect 2426 28340 2514 28503
rect 96 28324 2514 28340
rect 96 28278 250 28324
rect 2362 28278 2514 28324
rect 96 28256 2514 28278
rect 96 28176 184 28256
rect 96 16994 116 28176
rect 166 16994 184 28176
rect 96 16880 184 16994
rect 2426 28174 2514 28256
rect 2426 16992 2440 28174
rect 2490 16992 2514 28174
rect 2426 16880 2514 16992
rect 94 16844 2514 16880
rect 94 16796 210 16844
rect 2428 16796 2514 16844
rect 94 16782 2514 16796
rect 9449 28470 9511 28503
rect 9545 28470 9567 28531
rect 117 10632 257 11300
rect 2297 11280 2445 11302
rect 121 304 255 10632
rect 2297 342 2449 11280
rect 121 298 273 304
rect 123 292 273 298
rect 2297 292 2451 342
rect -249 -153 -229 -86
rect -195 -139 -131 -86
rect 9449 -110 9500 28470
rect 9552 -110 9567 28470
rect 9449 -139 9511 -110
rect -195 -153 9511 -139
rect 9545 -153 9567 -110
rect -249 -170 9567 -153
rect -249 -179 -136 -170
rect 9468 -179 9567 -170
rect -249 -213 -169 -179
rect 9485 -213 9567 -179
rect -249 -222 -136 -213
rect 9468 -222 9567 -213
rect -249 -257 9567 -222
<< viali >>
rect -148 28591 9456 28602
rect -148 28557 9456 28591
rect -148 28550 9456 28557
rect -238 -86 -229 28494
rect -229 -86 -195 28494
rect -195 -86 -186 28494
rect 250 28278 2362 28324
rect 116 16994 166 28176
rect 2440 16992 2490 28174
rect 210 16796 2428 16844
rect 9500 -110 9511 28470
rect 9511 -110 9545 28470
rect 9545 -110 9552 28470
rect -136 -179 9468 -170
rect -136 -213 9468 -179
rect -136 -222 9468 -213
<< metal1 >>
rect -249 28602 9567 28621
rect -249 28550 -148 28602
rect 9456 28550 9567 28602
rect -249 28503 9567 28550
rect -249 28494 -131 28503
rect -249 -86 -238 28494
rect -186 25235 -131 28494
rect 96 28340 184 28503
rect 2426 28340 2514 28503
rect 96 28324 2514 28340
rect 96 28278 250 28324
rect 2362 28278 2514 28324
rect 96 28256 2514 28278
rect 96 28176 184 28256
rect 96 25235 116 28176
rect -186 23202 116 25235
rect -186 5650 -131 23202
rect 96 16994 116 23202
rect 166 25235 184 28176
rect 2426 28174 2514 28256
rect 166 25232 276 25235
rect 166 23206 267 25232
rect 2341 23206 2351 25232
rect 166 23202 276 23206
rect 166 16994 184 23202
rect 96 16862 184 16994
rect 293 16928 303 17048
rect 2301 16928 2311 17048
rect 2426 16992 2440 28174
rect 2490 16992 2514 28174
rect 9449 28470 9567 28503
rect 3343 21278 3349 21386
rect 3457 21278 3463 21386
rect 2426 16862 2514 16992
rect 94 16844 2514 16862
rect 94 16796 210 16844
rect 2428 16796 2514 16844
rect 94 16782 2514 16796
rect 2778 15727 2968 18974
rect 2778 15537 3366 15727
rect 1 12929 103 15196
rect 3176 13773 3366 15537
rect 3176 13583 3660 13773
rect 4349 13604 4817 13764
rect 4657 12132 4817 13604
rect 3929 11972 4817 12132
rect 3929 11956 4089 11972
rect 2775 11796 4089 11956
rect 275 11346 285 11440
rect 2285 11346 2295 11440
rect 2775 9236 2935 11796
rect 3343 6934 3349 7042
rect 3457 6934 3463 7042
rect 229 5650 239 5652
rect -186 3682 239 5650
rect -186 -86 -131 3682
rect 229 3680 239 3682
rect 2335 3680 2345 5652
rect -249 -139 -131 -86
rect 9449 -110 9500 28470
rect 9552 -110 9567 28470
rect 9449 -139 9567 -110
rect -249 -170 9567 -139
rect -249 -222 -136 -170
rect 9468 -222 9567 -170
rect -249 -257 9567 -222
<< via1 >>
rect 267 23206 2341 25232
rect 303 16928 2301 17048
rect 3349 21278 3457 21386
rect 285 11346 2285 11440
rect 3349 6934 3457 7042
rect 239 3680 2335 5652
<< metal2 >>
rect 267 25232 2341 25242
rect 267 23196 2341 23206
rect 3349 21386 3457 21392
rect 3340 21278 3349 21386
rect 3457 21278 3466 21386
rect 3349 21272 3457 21278
rect 299 17048 5021 17468
rect 299 16928 303 17048
rect 2301 16928 5021 17048
rect 299 16884 5021 16928
rect 2546 16057 2610 16091
rect 2546 16056 2721 16057
rect 2546 15975 2831 16056
rect 2546 15971 2610 15975
rect 2720 15972 2831 15975
rect 2720 15958 5910 15972
rect 2720 15802 5536 15958
rect 5896 15917 5910 15958
rect 5896 15835 5913 15917
rect 5896 15802 5910 15835
rect 973 15701 982 15799
rect 1080 15701 1089 15799
rect 2124 15789 2222 15798
rect 2720 15786 5910 15802
rect 2124 15682 2222 15691
rect 3570 12536 3834 12576
rect 3095 12412 4987 12536
rect 3095 12286 3219 12412
rect 3570 12406 3834 12412
rect 544 12161 684 12285
rect 2665 12162 3219 12286
rect 277 11440 3610 11540
rect 4863 11464 4987 12412
rect 277 11346 285 11440
rect 2285 11438 3610 11440
rect 2285 11346 5045 11438
rect 277 11152 5045 11346
rect 3192 11064 3618 11152
rect 3349 7042 3457 7048
rect 3340 6934 3349 7042
rect 3457 6934 3466 7042
rect 3349 6928 3457 6934
rect 239 5652 2335 5662
rect 239 3670 2335 3680
<< via2 >>
rect 267 23206 2341 25232
rect 3349 21278 3457 21386
rect 5536 15802 5896 15958
rect 982 15701 1080 15799
rect 2124 15691 2222 15789
rect 3349 6934 3457 7042
rect 239 3680 2335 5652
<< metal3 >>
rect 267 25237 5034 25260
rect 257 25232 5034 25237
rect 257 23206 267 25232
rect 2341 23206 5034 25232
rect 257 23201 2351 23206
rect 3344 21386 3462 21391
rect 2809 21278 3349 21386
rect 3457 21278 3462 21386
rect 2809 16150 2917 21278
rect 3344 21273 3462 21278
rect 5523 21216 6790 21378
rect 977 16042 2917 16150
rect 977 15799 1085 16042
rect 977 15701 982 15799
rect 1080 15701 1085 15799
rect 977 15688 1085 15701
rect 2119 15789 3155 15794
rect 2119 15691 2124 15789
rect 2222 15691 3155 15789
rect 2119 15686 3155 15691
rect 70 12509 2750 12589
rect 70 12329 360 12409
rect 3047 12006 3155 15686
rect 2811 11898 3155 12006
rect 3627 13332 5399 21104
rect 2811 7042 2919 11898
rect 3627 7610 3732 13332
rect 5256 7610 5399 13332
rect 5523 15958 5612 21216
rect 6670 15988 6790 21216
rect 7081 21092 8917 22848
rect 5523 15802 5536 15958
rect 5523 15192 5612 15802
rect 6670 15192 6797 15988
rect 5523 12414 6797 15192
rect 3627 7470 5399 7610
rect 3344 7042 3462 7047
rect 2811 6934 3349 7042
rect 3457 6934 3462 7042
rect 3344 6929 3462 6934
rect 229 5652 5034 5662
rect 229 3680 239 5652
rect 2335 3680 5034 5652
rect 7081 5518 8917 7274
rect 229 3676 5034 3680
rect 229 3675 2345 3676
<< via3 >>
rect 5156 21510 6670 26532
rect 3732 7610 5256 13332
rect 5612 15958 6670 21216
rect 5612 15802 5896 15958
rect 5896 15802 6670 15958
rect 5612 15192 6670 15802
<< metal4 >>
rect 71 28247 6798 28248
rect 71 26663 8519 28247
rect 71 26532 6798 26663
rect 71 21510 5156 26532
rect 6670 21510 6798 26532
rect 71 21216 6798 21510
rect 71 15192 5612 21216
rect 6670 15192 6798 21216
rect 71 15044 6798 15192
rect 7052 15053 8519 26663
rect 71 13332 6798 13464
rect 71 7610 3732 13332
rect 5256 7610 6798 13332
rect 71 1839 6798 7610
rect 7052 1839 8519 13450
rect 71 255 8519 1839
rect 71 254 6798 255
use audiodac_drv_latch  audiodac_drv_latch_0
timestamp 1721164599
transform 1 0 1480 0 1 39112
box 1834 -27002 3224 -22840
use audiodac_drv_lite_half  audiodac_drv_lite_half_0
timestamp 1721165872
transform 1 0 8677 0 1 35642
box -5906 -19828 176 -8926
use audiodac_drv_lite_half  audiodac_drv_lite_half_1
timestamp 1721165872
transform 1 0 8677 0 -1 -7276
box -5906 -19828 176 -8926
use audiodac_drv_ls  audiodac_drv_ls_0
timestamp 1724508986
transform 1 0 3778 0 1 31945
box -3728 -20005 -570 -15559
use sky130_fd_pr__pfet_g5v0d10v5_VDASXE  sky130_fd_pr__pfet_g5v0d10v5_VDASXE_0 paramcells
timestamp 1644523392
transform 1 0 1305 0 1 22589
box -1258 -5797 1258 5797
use sky130_fd_pr__pfet_g5v0d10v5_VDASXE  sky130_fd_pr__pfet_g5v0d10v5_VDASXE_1
timestamp 1644523392
transform 1 0 1285 0 1 5797
box -1258 -5797 1258 5797
<< labels >>
rlabel metal1 1 12929 103 15196 1 in_hi
port 6 n signal input
rlabel metal3 70 12329 360 12409 1 in_p
port 1 n signal input
rlabel metal3 70 12509 2750 12589 1 in_n
port 2 n signal input
rlabel metal3 7081 5518 8917 7274 1 out_p
port 3 n signal output
rlabel metal3 7081 21092 8917 22848 1 out_n
port 4 n signal output
flabel metal4 71 260 6798 2260 0 FreeSans 3200 0 0 0 vss
port 7 nsew
flabel metal4 71 26570 6798 28248 0 FreeSans 3200 0 0 0 vdd
port 8 nsew
<< properties >>
string MASKHINTS_HVI 3080 20450 4700 21550 3080 6820 4700 7920
<< end >>
